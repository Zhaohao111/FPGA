module color_selection(

    input key,



);



endmodule

