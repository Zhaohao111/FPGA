module gw_gao(
    \vga_driver_output[15] ,
    \vga_driver_output[14] ,
    \vga_driver_output[13] ,
    \vga_driver_output[12] ,
    \vga_driver_output[11] ,
    \vga_driver_output[10] ,
    \vga_driver_output[9] ,
    \vga_driver_output[8] ,
    \vga_driver_output[7] ,
    \vga_driver_output[6] ,
    \vga_driver_output[5] ,
    \vga_driver_output[4] ,
    \vga_driver_output[3] ,
    \vga_driver_output[2] ,
    \vga_driver_output[1] ,
    \vga_driver_output[0] ,
    \u_vga_driver/vga_en_1 ,
    \H[7] ,
    \H[6] ,
    \H[5] ,
    \H[4] ,
    \H[3] ,
    \H[2] ,
    \H[1] ,
    \H[0] ,
    \S[7] ,
    \S[6] ,
    \S[5] ,
    \S[4] ,
    \S[3] ,
    \S[2] ,
    \S[1] ,
    \S[0] ,
    \V[7] ,
    \V[6] ,
    \V[5] ,
    \V[4] ,
    \V[3] ,
    \V[2] ,
    \V[1] ,
    \rgb2hsv_top1/complete_s ,
    \rgb2hsv_top1/complete_h ,
    GM7123_sync_clk,
    tms_pad_i,
    tck_pad_i,
    tdi_pad_i,
    tdo_pad_o
);

input \vga_driver_output[15] ;
input \vga_driver_output[14] ;
input \vga_driver_output[13] ;
input \vga_driver_output[12] ;
input \vga_driver_output[11] ;
input \vga_driver_output[10] ;
input \vga_driver_output[9] ;
input \vga_driver_output[8] ;
input \vga_driver_output[7] ;
input \vga_driver_output[6] ;
input \vga_driver_output[5] ;
input \vga_driver_output[4] ;
input \vga_driver_output[3] ;
input \vga_driver_output[2] ;
input \vga_driver_output[1] ;
input \vga_driver_output[0] ;
input \u_vga_driver/vga_en_1 ;
input \H[7] ;
input \H[6] ;
input \H[5] ;
input \H[4] ;
input \H[3] ;
input \H[2] ;
input \H[1] ;
input \H[0] ;
input \S[7] ;
input \S[6] ;
input \S[5] ;
input \S[4] ;
input \S[3] ;
input \S[2] ;
input \S[1] ;
input \S[0] ;
input \V[7] ;
input \V[6] ;
input \V[5] ;
input \V[4] ;
input \V[3] ;
input \V[2] ;
input \V[1] ;
input \rgb2hsv_top1/complete_s ;
input \rgb2hsv_top1/complete_h ;
input GM7123_sync_clk;
input tms_pad_i;
input tck_pad_i;
input tdi_pad_i;
output tdo_pad_o;

wire \vga_driver_output[15] ;
wire \vga_driver_output[14] ;
wire \vga_driver_output[13] ;
wire \vga_driver_output[12] ;
wire \vga_driver_output[11] ;
wire \vga_driver_output[10] ;
wire \vga_driver_output[9] ;
wire \vga_driver_output[8] ;
wire \vga_driver_output[7] ;
wire \vga_driver_output[6] ;
wire \vga_driver_output[5] ;
wire \vga_driver_output[4] ;
wire \vga_driver_output[3] ;
wire \vga_driver_output[2] ;
wire \vga_driver_output[1] ;
wire \vga_driver_output[0] ;
wire \u_vga_driver/vga_en_1 ;
wire \H[7] ;
wire \H[6] ;
wire \H[5] ;
wire \H[4] ;
wire \H[3] ;
wire \H[2] ;
wire \H[1] ;
wire \H[0] ;
wire \S[7] ;
wire \S[6] ;
wire \S[5] ;
wire \S[4] ;
wire \S[3] ;
wire \S[2] ;
wire \S[1] ;
wire \S[0] ;
wire \V[7] ;
wire \V[6] ;
wire \V[5] ;
wire \V[4] ;
wire \V[3] ;
wire \V[2] ;
wire \V[1] ;
wire \rgb2hsv_top1/complete_s ;
wire \rgb2hsv_top1/complete_h ;
wire GM7123_sync_clk;
wire tms_pad_i;
wire tck_pad_i;
wire tdi_pad_i;
wire tdo_pad_o;
wire tms_i_c;
wire tck_i_c;
wire tdi_i_c;
wire tdo_o_c;
wire [9:0] control0;
wire gao_jtag_tck;
wire gao_jtag_reset;
wire run_test_idle_er1;
wire run_test_idle_er2;
wire shift_dr_capture_dr;
wire update_dr;
wire pause_dr;
wire enable_er1;
wire enable_er2;
wire gao_jtag_tdi;
wire tdo_er1;
wire tdo_er2;

IBUF tms_ibuf (
    .I(tms_pad_i),
    .O(tms_i_c)
);

IBUF tck_ibuf (
    .I(tck_pad_i),
    .O(tck_i_c)
);

IBUF tdi_ibuf (
    .I(tdi_pad_i),
    .O(tdi_i_c)
);

OBUF tdo_obuf (
    .I(tdo_o_c),
    .O(tdo_pad_o)
);

GW_JTAG  u_gw_jtag(
    .tms_pad_i(tms_i_c),
    .tck_pad_i(tck_i_c),
    .tdi_pad_i(tdi_i_c),
    .tdo_pad_o(tdo_o_c),
    .tck_o(gao_jtag_tck),
    .test_logic_reset_o(gao_jtag_reset),
    .run_test_idle_er1_o(run_test_idle_er1),
    .run_test_idle_er2_o(run_test_idle_er2),
    .shift_dr_capture_dr_o(shift_dr_capture_dr),
    .update_dr_o(update_dr),
    .pause_dr_o(pause_dr),
    .enable_er1_o(enable_er1),
    .enable_er2_o(enable_er2),
    .tdi_o(gao_jtag_tdi),
    .tdo_er1_i(tdo_er1),
    .tdo_er2_i(tdo_er2)
);

gw_con_top  u_icon_top(
    .tck_i(gao_jtag_tck),
    .tdi_i(gao_jtag_tdi),
    .tdo_o(tdo_er1),
    .rst_i(gao_jtag_reset),
    .control0(control0[9:0]),
    .enable_i(enable_er1),
    .shift_dr_capture_dr_i(shift_dr_capture_dr),
    .update_dr_i(update_dr)
);

ao_top_0  u_la0_top(
    .control(control0[9:0]),
    .trig0_i({\rgb2hsv_top1/complete_s ,\rgb2hsv_top1/complete_h }),
    .trig1_i({\vga_driver_output[15] ,\vga_driver_output[14] ,\vga_driver_output[13] ,\vga_driver_output[12] ,\vga_driver_output[11] ,\vga_driver_output[10] ,\vga_driver_output[9] ,\vga_driver_output[8] ,\vga_driver_output[7] ,\vga_driver_output[6] ,\vga_driver_output[5] ,\vga_driver_output[4] ,\vga_driver_output[3] ,\vga_driver_output[2] ,\vga_driver_output[1] ,\vga_driver_output[0] ,\u_vga_driver/vga_en_1 }),
    .trig2_i({\H[7] ,\H[6] ,\H[5] ,\H[4] ,\H[3] ,\H[2] ,\H[1] ,\H[0] ,\S[7] ,\S[6] ,\S[5] ,\S[4] ,\S[3] ,\S[2] ,\S[1] ,\S[0] ,\V[7] ,\V[6] ,\V[5] ,\V[4] ,\V[3] ,\V[2] ,\V[1] }),
    .data_i({\vga_driver_output[15] ,\vga_driver_output[14] ,\vga_driver_output[13] ,\vga_driver_output[12] ,\vga_driver_output[11] ,\vga_driver_output[10] ,\vga_driver_output[9] ,\vga_driver_output[8] ,\vga_driver_output[7] ,\vga_driver_output[6] ,\vga_driver_output[5] ,\vga_driver_output[4] ,\vga_driver_output[3] ,\vga_driver_output[2] ,\vga_driver_output[1] ,\vga_driver_output[0] ,\u_vga_driver/vga_en_1 ,\H[7] ,\H[6] ,\H[5] ,\H[4] ,\H[3] ,\H[2] ,\H[1] ,\H[0] ,\S[7] ,\S[6] ,\S[5] ,\S[4] ,\S[3] ,\S[2] ,\S[1] ,\S[0] ,\V[7] ,\V[6] ,\V[5] ,\V[4] ,\V[3] ,\V[2] ,\V[1] ,\rgb2hsv_top1/complete_s ,\rgb2hsv_top1/complete_h }),
    .clk_i(GM7123_sync_clk)
);

endmodule
//
// Written by Synplify Pro 
// Product Version "P-2019.03G-Beta4"
// Program "Synplify Pro", Mapper "mapgw, Build 1429R"
// Fri Nov 22 12:58:56 2019
//
// Source file index table:
// Object locations will have the form <file>:<line>
// file 0 "\d:\gowin\gowin_v1.9.2beta\synplifypro\lib\generic\gw2a.v "
// file 1 "\d:\gowin\gowin_v1.9.2beta\synplifypro\lib\vlog\hypermods.v "
// file 2 "\d:\gowin\gowin_v1.9.2beta\synplifypro\lib\vlog\umr_capim.v "
// file 3 "\d:\gowin\gowin_v1.9.2beta\synplifypro\lib\vlog\scemi_objects.v "
// file 4 "\d:\gowin\gowin_v1.9.2beta\synplifypro\lib\vlog\scemi_pipes.svh "
// file 5 "\c:\users\22144\desktop\gowin_fpga\project\04_ov5640_vga\temp\gao\ao_control\gw_con_parameter.v "
// file 6 "\c:\users\22144\desktop\gowin_fpga\project\04_ov5640_vga\temp\gao\ao_control\gw_con_top_define.v "
// file 7 "\d:\gowin\gowin_v1.9.2beta\ide\data\ipcores\gao\gw_con\gw_con_top.v "
// file 8 "\d:\gowin\gowin_v1.9.2beta\synplifypro\lib\nlconst.dat "

`timescale 100 ps/100 ps
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="default"
`pragma protect author_info="default"
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
nGQjNTRggZWOT6sWc6oyraDUFLfWAO/HbLF6wXbCqXPNp9WCDJpv1rHVczOIVgncR/b0+UeSwebZ
OxlPzCeuO1qPl8FPTKiUyycPd+J0aSTr5vl+//g43DlAnrAZWpp+9NwkyX7Tl4KQV38q+/ZFnqAd
fKrxDpwkhDu4v9GmdKTtVryneeZJtk+qfqQLeux8ui4DI7WokBCiLCcnunBZc7zPDJ4RNHhhj/d6
kphLiA+2e7BZhQi3+S17OFvZZeAZqB9QHyWn8tsgCw/p96pTPtatJ/h1TGMYgxgbBmCeWweLMmye
bCwg5pbhghYptD2zVIQFJWuiylXMfypQ3ZpFdA==

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="GoWin"
`pragma protect key_keyname="GoWin2016"
`pragma protect key_method="rsa"
`pragma protect key_block
x5gHfLwQ9h6IkqXYFQsKYOoMTbgAOviKZwc0Vf339pYT772gCzJCT3UDF+YsUsYbK+Pq7BKRT6Uf
HBulNYuf7y+Ku9k8h5gb4vT0dUa4DG8OSdHb7R0AC/h0AeBTlns2hBJ4OSQGxyyNBp2s9HonSdOM
8ZWZFAphVVtPxikUpfU8q9qzyHTb9jMLF3VfqHt1hy3qcsmu5t+UPmv9c2zjTl4NXRMUl5483dXo
fMq4baFS/ju/wiHFuRhteazMg0mM6BfGhtM2aDlFaVzlnFbwItgar6Mu4Fk1u80ynR+wqXfj4ur2
96zU62Pm3UBbG8dYUGOAgfAhYDkhAs6USGbytQ==

`pragma protect data_keyowner="default-ip-vendor"
`pragma protect data_keyname="default-ip-key"
`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=7104)
`pragma protect data_block
S64wz9lq30aLaC+kL/X10osfDUSymmrQf6hdQCYuLnmlW6w0Fzin4aO0g/WUobnGsoCOY7+vwaK7
shINCGen4o92p7HrSWBdN+5Baowett5dwKHQqJmKXDf8kRu2EUM6L5usvI7gmjwb0Oqr0AOxGdMA
IEt240OIHMHC5+4DWcK1R5uW4oisAZTZ0NJomTQDaMYTf0vbCXRvBfHpZ4l5DtYYykQ+1wrCdaX8
sSH+7Kja8QmLHvKxnpa8f5JIgVG/ucAiaLjJCwWMxb9Jgg651lo4it+/5Tpuo5y2qsnz4H1JMNUn
Uj2Wb4mlOEYAAuxfOQgISpA8CPBcEc7sbHGRaiqACMoKpmzuzNxNUD8P5cv6ovUqQfJUioqy8RZU
ncsdMPHyh5mNATv+rgnC5o/KV93EFFByE293XvqXEYEjt9+B0tjML3MngPfTex/cJ2bRYI1Y29hm
XTL62PjJKbMzmK9NpFeIkHzsZDbc2u2z/BIavl6tVtDLm+SAcnppavWyK/5wQreqZ2yB53u9z2o8
LprLjQ9sr4VB4syjJwQmDoIF3R2IbM/QcfbvefBq4dq5wIAzfUOIsG7ArZLpKq5bpD2Zb8A9OHiX
uvKXXGCAt2zRRcVLod4NupUa6X2EHnU26zdjJmoMtd40HPn4cS1oNYsj8oDgnMRuf/Usf2EPCPzZ
zBwI1jWvbx/LDqAKeiJy5p6Z3ppYHfexLl4KVFJwvZN/UAIWIEdE4gMnasijR0V/X7zNIff2Z+mg
Vst3itLdrWLhIpU72gmh+FTfXmgP5G0QzeUXu+8N1eSeRol7/A0ii/TmT6olTEgp5qz99PEILD9D
dwbTqx6rbR/vbvZYn5A6MKVaJHf1Cf2AGsVHwSde1kyO3hEKtQ4r9nRWUIdDLZuN0jDbKAOGjSOj
cKQrNjYtn3fCdAE+vAydqBHJo0aNdCmOVR4Q2pRU6nYrm/btQlG2q7hLFtC/KPp2DUkDmxN8r+5B
jtXBUi4kv0tFiBkb0PSxuTRWBbmxgMHvu2TByRH6BUq6yGS45JSdbjpP0iYwguTga9uQlQJseJvN
j15bPLNnu23qzXFj4YABLhVMn3u2NXCFJtuYMqFQMW1J4orX1gR/oDz9x64hSD6+sdyOMqp9gEDe
0WZRRJAd6GzrepdeVLDl8wkUL5q2LruU+iqjEWV6S9w6E/+nxR01/BtxYLYurB06WOIux2dQ288m
+GGE3sZDqGx+4Z8RhX1zXr+jWRREuhScq0o8HakXzrQJ5d6LY3XsmvevNbnVF62XHGOq0jtREcXU
H1rGoR5lC3ijAvpx7b8Nk6N9VmI+ia0y17PcS32wivatHlatOvDz21513YSpkq/Yw2A6uJRl8KVH
Jj+kLgnAtJuMsFxxnHHDEd0DwbhpHYNlklIcez4hcNHHcW8UY+129G8pPPfxT0aJwrvc8xdF3FO5
zGC7rZuAhq3x1cJ/zlTFsepDtjwvqoqUCODzgXBkdDzWftJn68ittbbm+zbQzXZHy39+5j/0bQGq
xrYRoc7uHFk9KdSbpbDJdvad2clSy0ty9w4csPYjbsz+kkb94vouUIdy2WpnMkdbST/cPwsGLpfj
udJD5z0gsk2qDLqeePnl3U/C9moYz+Cw5pa2tiYU0V8BmX7+oShtCNHaGx/694KY617H2GQzy3oA
m7axRdZFb0Wf5dz0Nx2TmDvYGlw8284EwrgIzrOmqP0aBAPXESpUujnN+olGWShGRd5EtgOyQLgI
HhCppZtOjMPSKULg1NinMUMFPFZIn3dNlRGv2wFaiFFWDgFJnKxRNHujBhtdwAf3yifrXHjvjlq+
rdBW/36IfXTsD2Hk9yW8sCyFEJ8thBI9kX8v9IynnWfRY77pExP+MXu6n1mMsAGI5+NMIIvtD3/I
8xOHQ4Fm3nw61qa/ENEbZE2xLwnNBdbKhRkOJ5E61hofSr+tdUO7JXbd6HEDKhyQgNHJRVAlCaZg
nxVNBSyNe05LUxwkXsArTwvBn8XteTvnwreP7Rvd46oUPX9at5gkj45CfbJkoid5ejxoP7oRA8pc
b+LtAJCrMLquvMjrcRKEjqw+yyUwIcTu2KqmtaORXZbFfDMTQidCAL5iiZiQBMmtRO3/2JWSeO/z
yisWQmRAJxgLaoyfQTxLqqv183VR0dQI10GRQNDUNkuSEADQyOOj93ejJfRl7bMQft7oV6nVSCuQ
y4cjRGk4zWKW0i3x9RhGpv3MBr3PSrgrf0dmtM+SQAyshs8XMHzJevWf/0Y+78vbIDJJg1KwCgc5
uDOLVwDKf4yKpJU7loF9aKfWzRojoC/RpzyT9A68n5qc+QDWvPhUBWhrKN8weI5h0z8dGcwY+9z9
yED1Ockg4xGHaqcWGGWbPa5C1rZUCPgFkHsmyLX8W66yGl24nohnk0O/GNwCNhNzhVwQwtkawho2
o4AiWfYhdFKXouZ/racJoqYuoAV/t9cIMNZEG2q8vvHIXNf6/NB3QDyyNrxBmJYSwEABPH7rCvDI
rDzMLY7dGRZ1CgyuP2Ge2RY28vqO1sN05e4EbXxxz2GQTnvAf62+oTQg4B3cMKNkFUzO4xLyV4M4
A3r8mmGj/Kw5MHLbs8dl44f+P9vU/+N7IiQWRgPdfhrNIPYmrRRw0o3UEl5GQMa7ersm2H20+i3Y
FLw9medsYw903pVmzIBH2R1YUdNrYOquqVdI3cEjOHbVLruEmC9CEP6s8mRyi9ixwNK1ZGF7StYb
lYUvkpMh/FbEOutMh2dAYwuCQaKcUtQmP3d/SMDOgrDKXiJKqE6tzq7W5TDy5HWT/Y43/TdUF8BK
0jJX/krAu+lIqq+KfAkrBVy1aZR7TVrpuJptvSWUogS/ZKOQecBI+DScbiM3p7ZHod5X9Hlt+on0
Eix/WyX6Xh7Qr5AqZcNwvF6rTmcIBKjZv6j+y2Flnb7VMqDsTB8bAOoBRPnWW7yEWyy4GXrxoX8F
Pj4hlK/sGSmfTI1ioE/HOfBGFUrMTCaxpq3uOcMxBQeeNoZJzL1HfxDFntp0z1s/Rv/KJcGluUaU
LRAaH/I5r9XgOinwSRcjpBrxjS+uiwZXJu1JuCQz+pQcsbsP1hc1ZM12XHKr/G9/xkPgzCiMVkLk
E0wlaFyCxuwgxb889oZCDYq+huWYcNbgMGyi0aW+QYuE8Ha9YlNJf3A3XJxk8tTaxhWqXNp4THVn
ZU7UM9mZwAvK6ef4+/UugG5R0gLQMPPSa4+TeXQDgSYeCOWKs8fwhKrEpzgFgoPv1e20fd7MS/bU
Op1AIbsXYQcxcPvkx9+QPszLjD2V5z1vmt91ndI0sgzflNwbUVdkhMwrBYowMnJKdCru7q6mqi/a
mCV3l5rBjDVHh0LiICc4jMrrSo6EiLhNwWFJWowZWTCkUNIZNUKegYjpBs7gmpuwndeGNxVfXCZn
iVlTRNTIfWj2fb8GIQ/mJDa7hzFxv/21KhESvnTDuaEjy9HaxR0+OljsYi6owDKtW/cj4ei5Khnn
kKXigqdMoPQnBBy5+Dlu8xs2AWSIQa1wUyoGqjBATErO6LXslghIbgq3y3ExZTY5kf7IKKLBmQaz
YxJh3X/LJLQkgk7ePJveOrVRNEA1BMm4TdqAFj4pBlAUeMcilNPhQ+gX38QGT480Pc2RFSWW1+ZN
oefjAnTTwBcZ8z5Yac/0qMttIH0mDph96GRuSx8VEpQ0hr5VAkTVoUohABBRUHcb9Ls90mRafwUA
lbI3mwbhRsCkcsDJB4jutp3wOCt0BVnc3b2+PBN7AjQRSASl93ofLhAxfVQ03l1nSibvSWe1+wbG
2dUJy5u2M55OD1N5tEIcI6o95cLbNOx36bQSpDSigg8keHtqgKYe+fFnQZUWWXohOI5mATn5hRPV
KiZfXbB31Oa5A3DDm+jb5C4+D6mSI2LLcQZe6yknElDChlD9GQhlBTqUAG8cGVwlMftOZ5E8BwPe
rkBZP4Ih+w5WxPnkeYmydhqWLnoSSI6HIFK+gkJzsuTlBOU93wYBBG6Umg67l3bAjI4Xib3N5jiB
ZbFxokxItCnNtf1FFaLK0+2KHPTAPbuhOE2o2IYQpnab8Zegs05TYPyRSf2/7WpTtkDdiF7ejKlc
sPA+xM8N6R6Yrwakae3dS+Mu2Y6OntbT4U51BJmslkUEf0mWTY96RF1BVKUL5SVRgCqHRAeMyHaz
qHvSApD1czKbgf4i6g3q68umeUXAJJLiegmNd+yLjbdIGrlofjvBhlw3n6umwbU2Sqxw0NQM8HQ5
K6XxvdnDQ1OBfko4XHIFhhkhse8agYli7HJ0cpOsC0vaeHoA+BTC0lAKOkOLLD9Q+wI5y2lOBRUI
R/+2kC8ndhlEWoROS1M+bMQ8AURisonhvfmHAt62wu6CSGlbYwkp1I3sUxtx9kMmPnGSe5NHe1Jr
wGSchJ1g/D0weviUf/8UAtojoJiQUi/eezHzww2DQfz5PvREUkVQC1Se72W8wF2L4ATqFFaua12b
wGFTzC1JLsaMMaPmL8v5S0d4vhhorHtY4uzrMjEeS8uzcjyssxaVOE/ZLklT7bX8DKdlmIhWRAKV
qHHvdKv7weZ9yTsxXKWZaUpg4MHP0v0gdGecJ8xkSageBrXGZp1pI47y6W0v7bc3EMyt7rV7D2nM
hwUGuqQhktdwoQiLapiHCtuLi1cKGeScbabmqW0gFXV5ooMTafetu2mHFAhx6q02YZAPQhfcosP/
gwCqIcK1YPBEyJ60SkW9/KGp/K4XCOuyqgbcI4RHUPXCHgI8cVy2pRTbCRMb2mi3xA/Z90FEU3Xj
uQrcGrPom8pyR5E+2+9LpynAldtSRq8Zcv5RDP9JX5UzC46Wz96g6N+mgtkn2HEf65hkGMeE4lHl
7QkSgTEPQU95gFeFdkSbRIzkbBuFoYeLSRg+C2NVZafssUKr+hmVdhlxpaBI8H/Pm8bhBdMuTDXe
baF4PjmAlt+jvXOW//65RpWxZIA7UMjfPM0qvzyqNa1pxutYSAlv2o1PcmRbP4FWJgREZrqHDODh
tH6WmdjzAX/aekH+OByWGjNbusM18D6S4LlsGX3TIzolLYTrISa2x6rD/dhMH42XZ3f4Euhx3p81
JBGaLYR0T6RDiPaxX6lS3M5S/iCG33e7TN4pN6sgdSsnC1dGZG+R0hxlKTJ8/uV4NNtzkPA/n3Zb
V/Ygx3XbsyC5jh+IHQvpMLdvbbZi3eiwvHwY5FHbhbBG5/UA8B1WTNIozV+Inb6mH6Ql6upBbU7n
1BfBMCH3b7kgLpqj8FycR6TbdsifLKegykv4rvvIUfrFos4NRkDaZigtCaiIZnVXVpTO1pWb4zif
EgNlCkNstuHrqcoEPD3crhgsmeH6Xf/rz8L/q1j9Kgqpq9qPUwUmttjr3ADtq4sTp8OgyDp2JaY4
6vYD3iIlvsrZsntzpWMm6c9TPsd5cTVpBnUWd7aB7v0eMN8BEbrJcwZPQef53ogY0XqPYaEL+gko
csex+bKwfWUBCIa0CQFsVSMTJe9XfCiItiSDI5COuXus8rISVFLgwl9d8kiYz0wW4Uc5/jGhwGVX
zhQTdRp0cN9HA57fWmind5vjXwI0qe9yRK78v1upOq1Vmms4KMz/teObjCkPbX2B9HaUQiRhVt33
tNliZfjsVNVTY/oHA5nCz++NA1vN4U0qKQhI2MagqKVuWvCmdyqLP+lf8FTnYwrGXYeg4MOZ0T0T
WzhUhv2C/dNmk8N6/bBUkJuH+WXhb1pveUkLBM3M3YQIYKbjMZTNooiG8dvzTIWbZRipW0rfltGg
rxX98Xl4nw43GXLStEFK8zFBjSoYFqVRMrxgyT+1VKGR8kEYIam3L1ZeP2qWvw7+Yv6+8rFZzKeZ
fVjENVwZ+10eIBH9pHtOZtC8NMv9St1efR33q84L3UZ9YoN+brKClkspTGiw7xM6WMZxur4Xj5K7
3Ct95Si7wTDo7hrfsHA7EZhyCAu3CDJg30Yc8iHhD6oCXL5Jbn4cgi0JAiiIUmXu0lXra4o1OrJG
OEmhCcpHIaRtlsDuyhat8zQI33wGe7LmOThpLb65qT3WWK5DJVxnJb+BNALWwz0bNckMVcWjPjvZ
wbWRKCo3RJNQXFiYWGpDlujc/LoTckBnG42+9RtV5FteQdb3k2KWxs+EyDzmWuwJzt9tmff0eZZC
gktiPz3lhmWywZtI/GZY4E7D6zOo8f/Gou79Sll1LmKjrJoYerB7+BHDEkWr6bl+uR6LvuCO1NMh
8G/+IcsgDLbpZB5T0XfebVnp9EkfVSklT21oxBixgi3KSFOi9eWAJp3zXrTY4RlxpBXcMTr3gvlF
chOj9VsyNQAX9jp8eIZrx8UAZf0uBe5I9WVQ0cOGJDdwumtgdvmAwYyiHwzyGNZ0lUMkzKNMQtXA
2Gf0xVP0mkRcezCmiqoFTGu35veszVCnM+LYQe9Vf18LaD4Cv2ztI1+RjTTn996RNBHkUR0n1ZVR
/JOkPTQGZ2I7wRc+UDlZlZgbyPSSfBJJjoDBUuNGacDYSB5RMhrmKwpu4ej7ESSqnx9xiLQRCJ8k
mhlxgHN0L4RyNYLHfuQNU12gepUGGjy8CgrLxeV3SRDIRuWqMADgfDgLrypwBqPorM2sMs9ptX68
ktZFXcwxJdcqo7diINqZGmGrlEIfuh4cTGp2j0BMfMgzbeYUpfaMOC90U66LKoub+dp7aaBdyyzX
OSl858zl6Lw6wD+bMtiqGboc18KwIF7NyesiOte1SF1CjCbIawvMNlAO7ORmQ5RZyOUKgnkOiTBO
3vgakwZXogeXnYrZXjwAKHlPuWAmiiXRs1sBu+slXY6MDMQv5sp6AAd4wj5DD47Ekvqa49Im77Pl
NnCFOod0mtE0+999pgisGX3rlFq1CqsapTgnX4XvsCrYQmxZsdAdIbjiQxIWZZGwy6zAFPi/YY5+
l9MTHXZBO8G1+iJtEENsF/RXb2fdkDj/p/VhmljDFL5DsGk7Iuk+X8OrazniOoDPqXtFaPPSb8d7
o5CwXbtQMmuthC+kjoomZmrJ7SmFneiw9p39ckPoZA2RqgYsWYTMD0wcwAsTHe8T32VGjAxHXb4w
vTIAVNH5wpxDKNOAodjFMSwz3qBcghDJwctosIPna1U3oU6paurBSDH1fPESGHShTsuCDPkNt/3A
ymgFnsOCYBzu6zuo/jECemOIMVLykEINTED/91fxnmmgmX0J0flYvVtq4MNZ7qWX/Wo5ssrMIMkz
+US0P2+t56X9yc9EsClGzRzNJdSAzFM6c2jZIz+p/VjrgKuyT0lhQPWEw9G2WUpB4xTtPhTsjQ6v
mG8o48RabcM9zOjLqYSQR87B9BHH2pD9pf5QtXTDjkGO/b6++aycn4oNCN+v+vrgGJAEHC2N13cW
RRh+i/1eIU5DUwBhFf5WegUCuhV5e1aNoLzmgAGOTf1evg5y7IJfTgg0FsnHXgMwBEYgCtiAEjLe
0+Fs1Yd0yMMl4q3DKH7wVIpZQBeYYVM+ENr8w9U8jS8N6q0JPGSbCNA3GQaqtZvsL4+RiJrXe3xr
vUIoMnxkHHR+ix3y/23R8hvVvhnvOnx/0YIB0fBy/ema0AnH+iBSjFaYLM7vuJvyCr4Q769jzT5q
u7RGBNQo8mXXoFmEe/suMcTSbeSuK/hwYB12bAyIDoaLToVOhHryyR514+pQCMz5KgS66TV9D3oi
a/3e6C0Og1t4KWg6it+TGLGw8RGJPh0MXoqR7y01no2Rpjs7MzlLH3E3IYZambc9YpdbtDCasv8W
Q5wKK2d9xr7MAU9XOTwscE4Xv9d6cr/bfirH7Lvjg2LWz6KWEu/UAn0YQZ+V/J4VsTn/bVrk/eaX
PZpSsFSesf7JBcYVGbKbmSTCH9iYA3dW//LvyPXuTz5V3686tABQqe521AR3OcVGr/2VHkbt1upz
PvROv6o6kNCj7NZTUGGkn4ZIjnqqhPuDPqHlVtHGN3t0V02WlcB9gqiVB7Z2sGteiBHKp/yEXja4
WbAWTDyJ7DqA36BuJwDo3vAQFDA8/dAvepjqYD5r5VqbJqudRyjsHuOLEKbdtJGZm5zWvGYYoNw0
ARqR4aiIMMSp6nIJUdiKc0lWZuie+ubOIBGZoX6OjWbm6NGTODFAD61hWGFgoR9yL7yhLuMtcrGg
1TKst12FTuVTDpT519TrwCAavJu5jLB6vVooDxUWfZRhgJOub7NYxx2A4aj95j5s8TuFqqdLPP0T
H41qe26XL2EUnRsQDXFX/JkHH/mNpXkNxNqJz/c7h08UTGn0tsEMypIkGYBirhZWkRC6YBrKAjzJ
NkVXRmNFKCPFwh7DsIYwq0hUjS6fd5KB4Sh0Go2a7t9nBhMVMr5R9QHyQr/CGMKLzvgpaxXTpHR0
mTkHjJNAeWzNVdYzTWG3sLqhC/9dFOfU6F3FLuN3WlsEkpyv1vPQ9iGl3MND2k5O3dPIxobPRmf3
o0T1oRw3gEQ1Kj8777jZO9I8Uny3h5KOv7pbKlOWeCjWb6MJ6N4Ct0TDBq++Skyv6YJipDIhJKqa
pL9IgvVUPM9ZtveUpCFTSnLh9WPRuJOTkQoYQkSpyPQuk0z06SOUgBU0Oasif2RC0ZOhOUlalUQ8
iWlh08Dv79eNGZIHJ2wstW67cX6d2mOR1u8UerxZXwuOWv9t/tKoUYlGruZ3JQ1LwWVlk4y2K7/E
cXY9I9YCQPJrMV7+Us2RifXM900SRft/vmFecRAQ2L1Fw9cy3hd7YRBcUpf7fL5s3i0a11xQQxXB
fKiiV+Dg9Xj3a7HX/u0bcnQ2VDgemdvOJMw2cNl/Q5S6zTYjGpvaHwFCd/46YWACiRCG/5cKoN/N
ueBzxbkXfVAkf9VJNTy85ep1a+NzjfuaU58ahtvTO9miRK2ZbucCsOeak61+6CIbB2es45bLzRml
6xUZSEsRZDN3t+uvmw/ujPADTmMzltXFpRqu1MmSaudaOK2aDXAZJj4/t1SdaNwAi4rMr64MWCvM
8GSpZVXHAaQ9MRoomQALFHzCNXBftQALac4Vm154Rr9JdfpO+C2zRAS2zrv0jBukrxc+kjOwKyJ7
oAKfYroPTvkgcIknimdNFqohPzHvcSroA3qsC5aJ7jnQEYtqbko+0p+U6cC1i/x7G72SPOr2cWep
jMkU1vNJv7a30OSBx4zak5x6FN78jTeGb4CUaxVMBVHzpYdqllvYP+7PDZeZ8IJcJb9VHzWWL+Vy
SvQBtEM4uwrUSG6Bo8Ecj3HBEktuN33NYSeSPXzzuMySZdAALD6Es2xXigIVqPCQceUDCVOe3BlK
WHF5B9WHHOL1SmhGO2VBaGYunZCbeQdtI5p0jnTVH8yXQHq4WzNk/v+igL4NWTOOs4Mp/prj+wkE
BCttwh96l3EqP2y27GcHnn6z4FYKMueLuhDDh4vSVAReMFkyObjkr958tFwKukAg05mM3Pgh/LmX
3PzsF4PQXOQizNvIyNLkHZ3B6iWi8rtPs4KQKEu5ZOsbQC+9
`pragma protect end_protected
//
// Written by Synplify Pro 
// Product Version "P-2019.03G-Beta4"
// Program "Synplify Pro", Mapper "mapgw, Build 1429R"
// Fri Nov 22 12:59:31 2019
//
// Source file index table:
// Object locations will have the form <file>:<line>
// file 0 "\d:\gowin\gowin_v1.9.2beta\synplifypro\lib\generic\gw2a.v "
// file 1 "\d:\gowin\gowin_v1.9.2beta\synplifypro\lib\vlog\hypermods.v "
// file 2 "\d:\gowin\gowin_v1.9.2beta\synplifypro\lib\vlog\umr_capim.v "
// file 3 "\d:\gowin\gowin_v1.9.2beta\synplifypro\lib\vlog\scemi_objects.v "
// file 4 "\d:\gowin\gowin_v1.9.2beta\synplifypro\lib\vlog\scemi_pipes.svh "
// file 5 "\c:\users\22144\desktop\gowin_fpga\project\04_ov5640_vga\temp\gao\ao_0\gw_ao_parameter.v "
// file 6 "\c:\users\22144\desktop\gowin_fpga\project\04_ov5640_vga\temp\gao\ao_0\gw_ao_top_define.v "
// file 7 "\c:\users\22144\desktop\gowin_fpga\project\04_ov5640_vga\temp\gao\ao_0\gw_ao_expression.v "
// file 8 "\d:\gowin\gowin_v1.9.2beta\ide\data\ipcores\gao\gw_ao_0\gw_ao_crc32.v "
// file 9 "\d:\gowin\gowin_v1.9.2beta\ide\data\ipcores\gao\gw_ao_0\gw_ao_define.v "
// file 10 "\d:\gowin\gowin_v1.9.2beta\ide\data\ipcores\gao\gw_ao_0\gw_ao_match.v "
// file 11 "\d:\gowin\gowin_v1.9.2beta\ide\data\ipcores\gao\gw_ao_0\gw_ao_mem_ctrl.v "
// file 12 "\d:\gowin\gowin_v1.9.2beta\ide\data\ipcores\gao\gw_ao_0\gw_ao_top.v "
// file 13 "\d:\gowin\gowin_v1.9.2beta\synplifypro\lib\nlconst.dat "

`timescale 100 ps/100 ps
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="default"
`pragma protect author_info="default"
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
DI4rXVSqQQakdxUiFbNMpUcFqLtxiH/v9VC2fotO6RT5oJx4ujfd+d8ntglwi9SznfUhuCDdANfH
XYMgV7tqilOQ2ZawjyjFzCrZ5SPXrGgsruT0nRljnPbi6qkiFtugOcQTRLawx9T7//cBM+KloXTA
NW5UEesUVY6XIevfIUZGJ1ure5Ny3juAG8DwrfgVKoVsVbpFHGqkn14/CuCrPfgd3cNIeMnz2tdU
fIIQcJuw7/y7oxsPIHnSNjduB2VlABUbTul3/U+MLlIz6QrQXnGGd0gsk0VzmjNw5t92AUKNXFJQ
KgZfLCLpjgQ/ZbGsMSNTxIFdLQdlxHMJmC0vaQ==

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="GoWin"
`pragma protect key_keyname="GoWin2016"
`pragma protect key_method="rsa"
`pragma protect key_block
BJq830S/kOcQBA2JJ2q4S6I8jB9jjQ+2w4M1vD4Tqw23sKPDOhifxjr0/o3W8kskkjrPH5ExmJnx
4+Ax8NsC3/y94RfnMYtaR48dVDd/uZPC+H97z8xQbMlRtAPIPBxmvbm2XF9esKwvNQk33qXslMT6
Af5S+VRtkbzP466p8XNJQwyztsU9oaM7FXV1jV3HosbJuRzcKVPEOmo4Dn/DOSxaP8rd5LPjoLqS
+itgiiOB0/sBM3oF4lMqNh90Lt7h7dN75Xc5z0AOiCtIi7ReGbnoPIxpLrTX3YY2f7/TaNJjwe2m
A2muDv33kmPJYj0Qn1mVE7WUxAUWY5au4KLJvA==

`pragma protect data_keyowner="default-ip-vendor"
`pragma protect data_keyname="default-ip-key"
`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=60832)
`pragma protect data_block
3l2m8UONmp/7H9fdVZbpxpmXcLOYUQ8E9OKnRpvBGbijcyKV2E6miLv/2ZQ1wwD3GuE5LklYVQEd
nav6lulUEdcSwDc2sj9bGjuo+OT3vo1ygV0LeWqkK8qUcZ66J388JcqXSTG017oCXYPU8yu2w7HX
UDTnd+Q64FViL0pQ7bWstAZ8nXO0jG3QHHLcfiSE+doD2LlJ7S53p0i7mg60ajc34nvE7wigXIhB
OKg9kKKIKAo3VgsUYkRHQX1oIFkU97dvx0cA+4TcbTju4+bP0kKwu9Tf7s5QENPkKGKl48VJpF08
7LnOP+Ck6lOpYvaOlY0GrWUHZPGiQBjY50BH9lhDksnwIX1hzNFCy+lW3T7O7Gx6otCzfzCfOSj/
F2gDMmPak2dDzNwfVN+k/5v6Iu62M23ZuzaL7cHrCsdhGA5T6jBorIRRY9bPI3sp/3Nd3mkmxqiI
CDt5AZvA6v6yq2aML6GF4DiewPTLUp2xICbNYkDEAdNmkIynRJMno19dOcr5MfKwkGlGFIFkO7jT
TmZvg8TyOiS2ckcbMwZXrHZupoRwq0SLyPnfcwE83fsUKKB77gUaLOelLlbpJzTiiIpNS+t1c1Uc
HrCbF0y1vSq7l6DUVVUyhH2843ohecL31ts5Zzj/WShXZPfORQ1Nk3VYM/un4bPPq65qgmzBmysS
wwgkvdEncvvps51AuEbFmiVZBpPNqCSxt4E7LXRobGEVX82RxI1qkEBtXfxAsy6K+0jLoTrizRTZ
dLcpNqF0jMfRmnugnETDE6QATLxd7JqYVITHdm6BTqZjsthGvatRuqb1Eoep9Yd9AF/o9RItbCG9
2MldE1Q9Zt/byyf61V1CLnZtClmClsXcTyZ6UGbIM5omFG3WgpRXGG6OSuOTqcaoejowux9qRxQS
XUFkQuybuKVvhHcveZ4ZOtok5yZpxpnllphgE5loNiJFn9PpcOazq6TpjvhnPTjRd7s1tcfmPGzB
Ww37Lr+0uu+N3a7r8d5QtKfxUz5nt8y5PcQwUMI5OGslaY/ZT5qVUR7HoeNaHy9Fdgp2LoGyjdZM
XNLjuukAs3ymQNISlLycfkwrAgyDvVtctMBTO6f74hSYUibo49o+bgLkGhwq0ixGiyne0txns7C4
RQd+cQocv2oqLm8njVSIv7NiQQ2AVh00YAZH/fDuDG+PsFlP97q1RRlSfhCXOWHV/PXrE8CqiXcK
/6psiaWgI8gVdw6vhuA2d38sZ6LGhZC7S3tysXBAmiO8WAJENm0Z7PVQgQXatpz10xW09dyv4LKz
tPU+PmmiLYghUqJsiAnni9NuNCaLZ2iuR54tUalTC+Ns3vsBMzJARnimw10T8UMuN7wlbEgaFIXE
nu0x85u9uD++pD6f2zZqHS5ngxu7w9o7NACPqu17NANhFmQcyioI2+19M1+kbIwH9OL0X2iKwnT5
C/ZjXldW/IibPYKld+umvq3iEREVjzCmm3ogs/cjRKbp6tWp4aWq9m3B/dQUl1xmNrpeDABFRzka
LF5lcae5DWNac789sRe4PnZGoUy5FLQXCPRdOnQOKhpSoCwtXE/NcOuRrfc8UqF8/qS9WEpnUanD
egOfXJeHdi1knB3eHXRTWLin63pknVcThUOjOehlIriRAjsTpKIx6GrcNHT4U/Ugm4HaCQOAu7A+
swWsoCyXp0CLOsH22EHX2R9GGuA5O8WCmBNofVSDfqLGmk0NmhCBqsSiaSFdWZy6O54vBUSDvC0M
7i9nS3NK3hge9wVo80Ups7g11HmwM/WgFaXT39v1MsT2Ebp/y6q/XrF1KeDdeXgQd+/KO54Hw8C4
aGL1dCewGhOfpoJHELXPQQR8GROn/WvZe4T1qdwhRSULBQJLvE7HgXTPbIOnJNqnixf7nui7EDhL
IrmoVw7z0F1zzZlT4CAs8/J8aO2XI+CUxxqH8OD8WZwlv2R8McR7VkVykUj/c6vpduIGKiTCUhXK
xGXLnMOreOLspfderZuh5YQdR9azhOip4MAQlY73qMPS1PQRiYzbsXEaZr3VGapXfU3bDO7LlAQZ
xLLdkdH9RKkS5TyT72lp4LuEbZTiNDYAMpn3gQ84PSxKyW+DwJTgByK6iVqePP7PfDHEtLre7Tyf
9TeatPWdCZ2FKgHnLPsY9LMcWQSfdZs8qP+Skg4/o3vpIQ88Qz8s02pYinWyJjCzn02kam1Z7hp2
HIgW22wPIq/xHHLK3pd5bw/gbg2czq78UYBwPmFtE9xXDGuDhsa0eTNq2YcnK5Rr4QThbiNT/Ja1
oHXDFM7FqIFA6yRmrLx+Fj89YVMJ445lrAeMbgPrYDYjRQcIG2fcZU/O01hYq6ZWjHj2/vNFpMi5
SjpIKOyFitjbleo6t4ltms04bEa9Jk9EZsTZFYjqHkSgJ4nv8Cn7W7gql91Y7zI1Edwy+8TE/Crd
PVIsbxEyftU4i2B8NiiV0ptzzMm2UZ0Y03q0nO+3psGpBPwecwOwmP1UbXtsD4LsABgEFmw8vmGY
Kam8HEf+n9FBa504t4AZwPpKw9diDM/25jhk1lCgl+vDjp/HsPRqpQOTvnWVHkSM0iKtecICIf+h
0sZ5htBMe/l9dlHg/H+plqlwmtOq9jM875Wcu4R+eif+4vbbjpeS1+HtZshZMsKs63pjpKUa2f00
NocUI3NGeVuWSgogcFTsk5geHwFDwsIudDGipRm9pALQBxqBoQin01/Vfyiaw/L8psxGzjQyZYM7
d0TFvuUAQI3g9O33pf+1hI1FYJK/slCYUh77xJTy67dQcHeboleiKY4AhRfs0gOlIo2JzkXeRaHm
9I7AKNvWpv/Ds+AOYdeSOHMEe06WutPHQZxZ0g+/jx4G4rSZ7Rgo0HliYvGwWmaNblyN3R1PVQ/M
IJ5UOd/+HBgVhI57UYqTWScPHRdraQLUcRViXiPMLo7qqjeCbFzf5IrWkJzwBz6BGsUaX9X1Tikr
N7jv8NE/hnuoakreT2lDiq2bJwrblV30ujpvpuSkcLZn+zg23qy/mZ2/mGaExz+oEzC6i1aRatTC
7u8uNFL1QftDHgPN+/ULTpK6b/EAd7rGOEMH9AhyIrK8tDGQp68gCR/zwd7tzrjwKJzj9Pw9M06i
QesMDizfhFZz3fXcZMkIEl5ZLyWBXEhTA5jY7r953MFYPq3iHwSVAZXhPNf7l8RwyOfcjw4uB+Tl
N1nj9tDy6TnCPxv+PapDBQs/XfWK9j1ICD9ey9xtyv5+c0oAOl7VJH/r6iInsXHkkfRP8G5iIJ2z
jIaKzO/yKnKuk7b/QoxpxYzyfPzmbc6x3iOmbr8Zq2r0FZGMzV8SfST5JKfIti3WuBqjTKCZNiQQ
gnoGw2bVTQvjjS/U0nqrFI5nfnBxXlBNS5xvHKE10s7ifmfs1fkjBsP7jQUhPX0wKSitOohI+s27
Lv2sibteQshwtbyFbfiUq2kfESafo+bdwRp9/g38a//2W/U8sSUWh/50rtMUem9t2iscMzLVK/jK
b00NdG/ZpB48+yxPkL0LXW9c39fIQR2HvS/8BonTUdFqcLDCJGcIhBH7xpe6rG72Y/pefIDurqXn
jpNQJmv1rvzV+gB4XUuJVn2vUyoGR0VVfZpI/oCP5TBDi+4iBYchIqCqUoYQGMB+U7uIN/F0mQH0
ylPXrPj3+bbbMRyYgxBfnnR5ihZ0oVYXpGxydDv5UaCYd32Agqy5q5f7gPUkwF4H8K0aGf91smy/
cMY59KJfEePrkLhWT6FMSaGPHUUXKxE9SzOaT1uPcGo8JQBpa5SYXtiUO2BdfNdkMgtYiVsiOiRZ
VAkbUVjW/3iAHbeE0lfqm/slrZuFCynnd1NnrUkArtP04LPSEL9SATnhXzVNmgsQ9WGX+2Hq5de2
cCzDlc5bNbDyQFCatqfUDAEFoLTMTtwFzp63hvM2/xSjSais2qmpkQ5e9CDOI/YJVz1NemrVj6AV
XMXoO0tHkl9qh7iE1foPEM4obJwv0hBtvtBg6MPFc1XhLlxhl1SUTKISiL2q+6FzqKOgLm6Ze3eV
UGYDhyJ0STDwuUh2Ndxje8Dcfp5iowb6ruOR2dr2H8OaFRPBVDaTpOFX9/YUuEmNTW8oi17QB0f4
LTV6QWHPW+09AtpTs/4X2bLHrILJaFjQSMP70dkevtJ1NnCLBu/4CppIZGKZDc6CD1JsFl2nMB96
419m1YUm2GQI8DKK7M2zFIskEZ+Me1hK/xc9c6ZRKQvEQ71mxuokoBywja0Yl0YYu2NjqqRPw0cu
L78/qEfbpViGiaGKl9/nZ2HZGhRB0+VxcH6oPWCfprqB6M63WTD9Xoc8zbFI+1YZdBFbsrEqGfmU
ZLJksbB/9PyQeoScFG5x+GMcZFO7kMjrSPR9y6HLYvLMS/cjzEweSIpV+KThoxztw7UHfGhV3Xky
0yTQnvGSC2Q/giQfdhVcPklNjJdFiTQ8Qe0DVxWHVvwpUkGQqpM7/4Iz8lcgjeke4+hJY2id6YMk
gOUOIFyLQV8NVkZ1VUoHfRIkMjIe+YKKA+ixB2axlhYKtKIm0S91TyY+CHR3jodkFzaWKFA03Chb
zePVn4acY4AfPvuaHM8JB77TnZbn9OnuNTV0zzRp539/SoGIs2+zlHQzt7lvoeuIj/weCQa93jAr
Aod09UZ4cdO4hsAB+Tlg1uycNMAe5bzMM1gFyPEwy8mAXRcOKpMlyu4kCWJ1rbbyDWddXnSRHqTO
RRjQl+WHi7e1f1nQsDrZb03vLIWcQn5mMz35yEWivWnrk+AV4Mtkzo8j2IeqGI3h8irL9S4E3oiY
T8WDt/EOMtnlUpjdcbvdutJx15scH8ID3sev/k1yOycnApxwrxEYTjcyWNzN8v0QfLI5DeM6Xfwq
a4It7v4biny/eyQ84iGSMS0Oi9nVJop90kSxKY//jFYGdyVijRWR+tRUZh4IPlhIYVpaBuYwFOgW
uLp6C6VY+pTcTKJiU97zXekLbmNCQNohXhJKmwkTyadXg1cBE5UFTDn7bpVTM9CVSC678eKdA680
zZ4U015SJzZdgXgPnMLJ9ZcNR7RzSJ1uH3ZkfBpVglprO2gm1XvKyL+dFAhiv/ViSi7Rw07A1GKB
ZIvQiUkVeS6fyBci9pU6mEHPwnm1UtyHX9jszMWYj52iOYSi21Q/M2+eYkquytI7qkZL6wx47gqR
9U76MJt2hnkwQTlhd+9WmlMJOcH2buDqI3slE26nXv2tW0Do9nDnsxEO/JsNR9bRBS6ECs/3U6hQ
4SqCGQrLCG4I7tOBatUZk0mtUx32Iq9RMUUcQ3kuaNavldOodCV5IbR4boxho8U2xjdcJ0Q1mRtp
XE68+H3iB4icbwpDWTtcyCP9FVxTLZqoMfc1gVRlZVNiHVuik6rl9ZlX9owK9t1Fg1as5mQJAseI
OEIZ8LkgR6BFmcLxSGAEfa7V52Rans5kJpweDFOxA11Vy2KdLIkiyENsYhjRInPpVZoEudbJK+9X
Sw3rxYqGiTIX6eCWoOitbM+YGDa33dME+GdQ1zwokCdEaKdAOrA8bDWkWDKxZMEoFde5YNP7j335
+Ztqa/j9GEBGnoMMzEVk4Btg390GqIOF5QyvgneRc0dZguxtK2XfTyPB0kfr7g6j5dlqpHvPozNX
mARX7rT+tvL2eJzmUSlto+kN7KE8L20W3WzWlt7I+f/M7pVgSYK9oaBlazsprKWBeGn4LBYDxRSL
KD8LrGnlysxYNdC0kDz5/iMiGI/8uSKtROOfyOCmXzTg2fJpai2655svyJt96EaayuxHT/BEhtnG
ouzrJEeZh37e7CSXiPtwvZw6IbgtEOmsqTypvmmzCE9zOR4+O7Hv9bG/cLzstazhBd0v9vtHuDIp
bMq71acipOF32u+wUQe6dJLg5LfdaYpgsnx3btwbOXWZf9ZK/2jFb7p6amko2LXKG5YbtG0CfPlD
zWok7YX8dBuFqrZ9qTbRfQV4LraZy/j5EE8bLx9N03dkwPYCAy2VEnMQhZSwrvjnXHUvsiOxLgsO
bDwvFTyIGdugWpYpG8bGwrK7OuJH7Z/HyaqPZoC31Wpaqu+QocW7lwp0XCbbOjNumuew/TxaeTBv
6Di6R71hgomA2walBX1QtmKoe3u+Dl0DXH2Cni0gTQ53z1SqFrktZoFl7cOt0vq6JdqMqHFeY7Zk
jGUFwD3ZCIZwKPugJVn10i6AVF9EhRXB7MGEZ5o5AzadryKzt2mX+QwjG/hjhG+67u448SvDyfIz
88ityQ1OF+2jYyoM6QNOIjeH2R4LErigjnJYoDOfBAio90o8Zwnycf9wtfJ/aZxWnttixf69tLHE
OYoo1pQ0Ygh6S6rQXFiHwwTwKSC/Y16XBwu0phFQE3OzwdYhr4Lt/V69SfaMwEIr1lhSIkJMdxWj
FFw06ezaLlVpqLuGoZE8y3OQuuJCsasSoFDAEheT1ndkwWTZhcOfocVD0PoONoAXUGWXYoDUaURd
fm5skvjt5YsqijFZ7iN3a4ItyQnzG2sHbg7nX+tS1JIz7tsFPUVjy+v1WcFkRG1N4IgZhy8JuEpI
J2L07wEGHZRLgDQbBNP3UwbLS9BtyzKWADXvkbaQmaR2vHMbV83L0JeTDjDzWymtyIX0WGlmbdRO
GAIsysK7ti1fH8wksI1bfWFbSZVbe8B4EiU7YVoANXWdLAC5Va1Oq4gpPdtMxR+SrxIfsj3PKGSQ
1yhadKH8JkjcnoGLxLTQiKJbof2Beunlx2iBAp+0tcWPy1HEAz6X0O6AO6fD1Y9PrFjQPE1kJ9ZL
WwN2/Vjbi57LwXo83jFYvSnqS1MeJ2QNR0slsleuj65Z3xDCuQVm7q7ddXDfNw/Z7jl9ROHgxGse
Rtey0OylhURCc18j03LITf18RsVM6A9IvNbnOXSd4I3FXrXpC++Am4py+mH422hy2hYR621qQvCh
3syOr8P7AH4F1daV7K9ZV+Oy1sjelojlD8hzIhiNWRaRy5Djf6HvRE4k+xkH3OaE1qEVJ4H/kZqF
EAov7SOt6SoprDp7ActBAKJ2BoQuNWZbwWWpIP7In5Vc0mE0ZjD7nkqBNZfvdCU85lv7fZOVQtVu
BzLOYLkvvL4YPQjrCIreoDcZbWaK5xo/+FQVlvqdjQSYjLzoFmCDWEuUdtPMkMJ8W7ZQkJUiHqxU
sajUcPiIKXry7c/y14se4JZUAljYqey0ilC81vsK2HqB1El8z8L71+Jgq/P1/qUKRGjiJ0ySaDZ7
oJK/VZ1Kure9gGdDa/eQjjZFiZC4w9nVX4CG9wYp7CcAr+TxqrCusbsY4bAxPoUnZidJ2zd1V6sC
cBOGXOFHZjaFyhJr0VgfvWtAiSS2WdJbHeMpcNGzxg/P7Lm1rDSFo8nDv4ah7Owr0crCVIm1X4TT
NtlGXSLuyOa+DyYeDmLSpTBFyACHNJ77X37ZFBLBCpxpiHlDk5iblMl/JoMhEFHlfCO3qD8rWeHO
d2uRV8l92duDfJK3Mmsp28RzNDtpfnOE2VIEphOmHfgVzPkUkxUF0G3l3qSUajS7QJoLzTdWSxs8
TugDNK29Zu0wVQAVk/bwLBO+KAv183e5rjpc3H5BXRkEgKFAn1vkqH/8+jbigCkTFfT/oC0ZMclg
7AoSXEbBAAiJqX6doGkz1A4JRvdVSEudwRLfrH7cozCuzntWFgJIqDZVRRMupfREF6BwmjahLblX
jlxas0YkCOYPmgkcNev4RBqCYBOhpIDf3nBSdH3BHAJpgejeW1DCmgDL4wnB2Oy9hd6ajrlEPAVi
/tGOuc96csrbuFjnz1TVdCn9hQfvqKQ+IWOpP01P6jI1Dqw0fezU1sQ0FDkJO+3eMbxPBW3F9IYx
OIDBJC6ciSKbkN8oNpgPV+EcD44AK+SAamNjtcl67o0Z/veg9pq9pM5yf0OF5mnB7IZP4dh9uAxe
27jEPvPB5TJqwOhE9ceQNfegaPx2nqznhqk55m7qeZCHvthCV5QIXCSqhDlTlCTkAZcxSGH1TLpl
d5cx47sD7Yrv3TlENT99F/vlYLFjhTCLwsuRcHZZStrXXA8tbUcCBCHNmj1ISCFtzacp3SCrPqQh
QiI0KXm81ZchE/iXMQrVdUfM3J2afnDjhA6y9D0mME4K0B6bc5V3DPzpMbsE9avxSfO4emTQ24ZW
wkC8ZYqThTK7lNpvku6Sn/MT76yMrqtwlpK2SE13FzadnxC2c3eZkSi+zi6tHuVugv+I4F7X/c6c
b3J3l5a0kO3BPoFO+WAcoKrwUfbq+siY1BEuC0vnNyJDImSlsRvrnDFrPbmGzyJrGPqEW4KUqlVm
uqbDwJWYqykw/aT0IORi3q6CIKR0v31auF0ed5IvJicwAWD6w8e2QwOQI6PdWlDgksMNrN0lQTqy
L9eg4mDGPLNjAWAIQmV6W+6V7qEI+8OB1bfOtKacD/52M6MhJe3JBd0qf/B89QPtTQeKoH7Y+JVv
q4YJwtf2CsrrSK1P2jFJUDMmJusLIbfgWNi+mZy7YWtsrPvkXyvChItLsPA3V3qaOrrJ3P6k4XxI
5l6HZ7UKDIdRaKZTD+aYWO+9LC5Dbj7koWgCiSPZSoF7TSbHMf7SRytaDBf972aY/0SZOSCasA8z
YFvXsmIjJXCGkc3rYVquPKQbj1iPTgrRbiAV5KQwHbdjRW4mOi4D8ZvztEarcgWaQpv/iarv0z7S
LW8yzfknvMi3JM2CiYZNRyWlgrCk4zFN6nonOkx+2Sc1dJnoCfeF33Q+4MxwG5Ow2jne618Upq3L
ijjge8qpJ+PBbOZZ7hBFirwWcXxOpIFv6hVLsqTZkbSff0eEpy/cKY/AIyEhq9nsyMC3vk9Dxs30
AbFk5ifAWQE76qFds0ibJSP3KM1VV5KhNJoFTjwC7nI8sgNdg94JzytQjZfK4+dwQV33wUki44Y0
A5GhnrI67JSDHfAitmk+A8rqWPD6Yng8L8SmFTUIO089zQR3RfPNQoVR1OD9lLsOczLVQeFA33Cb
popkZ3D60/zCBwW5JPV/t+Szicu6fRPwQ6oZ6hndUB1lQjlHpXxlU+4serJZFpTLp4JGnOp0zZr8
M659Ud1k6E5Q3k1rQsXm3b0zBMy8xn+8tcPJl5h+dIjwK+cxFNBzY/g89GuRLa0cB6m1lLzYgu7r
Igk1MM4Wulyi0dHVX/Bvz2tYpqc+6DXVv2vqaCEWaMvdfQ4vvOmZfncixLkzKy798OuPlfCM5rLH
oO2zLNxpLOEPVLL5D04sg43QZpYzCYncDYSRmFdtjYehgGSR48Vy92ocYQvD9fIz72FP3mEKVJQU
/ACQOeRm9VGXWQjldrkecULyhhOGe3/9t3/VQf1xw/zcK/zF2wZ1MOzGiFq7tDzKjuWbQLQF3fzW
p75FZLVkP4qMaxAEWMR5Z8UlZE+d1f69d3xilNEPGBlkOgQ+hr9ANoCOIxV99QyjJovWWvbwTdoY
WnGZbjS0yrM5q+07nXK52/qS63JS6hmU0Xr3XjMF+cJY8SdUnzEBfXkPNuu5u9hiP8rihkw49LJb
k4Ge/VRtrVT1FdNMnz3rw9WAIoCIaI35hxtfieqrO0cEFROpX7w3DMtn0XnMTuCNY8xdxS+EpArG
A+C9d1jqjj07OewPlwohK2P6bC1YR/8LW65Hm59eMbSXtNQ6nJT4xAsDDCFpkPBK39Pcm6sKFcwW
RQrHjv/qM6b3xGdSS7NEYI2O2h/nNxSHZSpXU8i2PfUW5nlTTD+JlqLz+DhrmKBX9/tz21CzPWNQ
BAGM5h1WecZR42tOn9qOV/F+4QZrnyedIFoJSGFHqYhmUGAXm/k4fCA2kQvrhV1+ocbPcQS930js
kpS4Am/+rAPDSd0cr/Swv5Ci3EtNqycU16HDqpm1rglaqbYH+Ev/J1sMwfjfiuLtN0vBhQA8vh7B
w4BW06s4kBYNEvG2Pk9ucIGZOJb6J/ge34dcVD4nngX/cd2fNp2pf3bfKgoWgEBV6ZdBKBlbdB2q
A2l0mPyw2ecoIc5nzC4M9YexyRPkSamCDu4lrxbFDG5ULg3TQjFgUpTGwukTYXYVB/k5kG62mXIi
ULQSZPycarsu0cWrB9D5blMFUWuMABrLNFSVqi7g5mAEaZFB6IBo8ay6lxnwS3gzpMRvrqRFhEav
/Uw/Gt2c+iDixgM9/qw5RUKE4VOOz9mgr5Re4wsc/VQJ/czpga6MBW1jjyOR5uF7EVgSX3w6FEW7
8DJ2Gjr6QceYZXR61pzq2rKYfzjVQyTrm4NRgPqql9Q5N07fak5dqgJLUdx17t5+26Vh4tnOQial
Zewfi/BUbTUX+J8s2PWOX4gpb4vpe4g3UlyUqvjNgktkxwfgVSodHyPDpwtl0GWUduD7LhQ8TUOM
mm08xFzL2KQ2qAEciKvMkAJvqkhAqDLoXmZlfaHF0hHLYDSpvnUpRXGBVHmLLj6xK/BVwlBX3UzN
XN8CQEWTr9YB8IV5U/GfvKF6N7bb57qssyucBQTsO4YykgeZMqXEkhCEAW+UFTLWxw3qxy9lM7js
uQZv4K2vJp4JN/CK4YlG7xTJZu4kdeH5N6Abadl+Qzp634pg4dwXqv+/9aHCBjuQGUf2OvtAxNZU
L2f2MYtGRUFbzA4JjVdY+A7lz6unQVtjyFbELNkKewjCrcctTlNM5p7GFalh0xQF4byV2LjxfI7O
odGrjN/ZHWmweF1ImT+dEGiewU27LJ/gcwORTxfsSeQnZZFQzfXtdCcv7cMQC8RKF5a3GMJIk1in
eHOJepN3ua14DmGe0VMaOPlFgJP6XtrwxKk7Qko0aOjC9sAdbrMieSN+e/csWiVM7Zom454u+otM
6D4IfCDA5qeIBSjiGPpNAC4ov2Ag1uGPmm0saGHGP4Pq031czaaADpWVGmcMEE5IHUli9PBubf6w
utXCRc2+wygK0YsW43iXLsoPDSkQD5WgwqB1k1LZge357F9HFOOeBz7823IDW6a8IXqMQGdDHf+b
seVMvAOiIoGivHl2b9Z9bpVdOsiHXXfITZkwOuZdofuO8lZap3zCHr+5vxYJHgFBSX5MQ0qjJ689
zmckmUCGjKpi7AU6mHlauo1p+sZAFcfJYLiF/dTo3onRZWSDR3jzNKmqo6Y9gm1pY4a3oOXZmURC
+fhWRS5mAALTXGKXKrBH/bn8icaxlA4LtHwuiBbxmt+FrF21fbzAvvfw5GAOLl3AVJ1qctwSlHEP
kv7a8kacoNCEX/hD6bxDuwUzWg9trvRy74pL4xFcWbKjT+EhR27Iudri5ZaDVYsj07fx5Bomf5Fk
VfWvaF6+dBVJZS7nfRhLPbjpZc3lcQe4eT8W9dqKf06Oygns6/4BHJX7PPvpN0tTuHBfGKjpiQVJ
2vKDOhT+8pOI3NBgC/P4BOKzKhMViK+QDbKsqkIMBh/Fg03c2GnqneYH2eWntuD5eH52uEC9wY5n
dyrpbJTYVxW4PG83B4xaTUsj3IRyG7rs83EletDXzcElK1mn2wfa5bSP5nzm2WBVfZw5ypxKaDmT
Guo2jnR1vsgfxIN3RrnfJuCC6Dn79FR3NjLWa/XIbm835vvFNIW/ItO4aGvwBX4mbw2N1eg2rX8N
sRR19F0QaaHmzC6yTd7cO2GcJkXIb6dvKmYVJUTVd76OTWxI/fc+38hX1GLq8ulua5VFHjv1Zr+h
mJv5i4Bbx1tEd2miHhPwGiDoRChUgr8gM4kQfKqwntwzjLbg6/ckrxY67c1TSbGyvfadNgNgYeoN
ftSjsSVfVYd1lnxZbcBia0Fpviln2w4UvpAbm2VkkFqDztQwXD6GdJFSErPgtEc/NoMaRUk2LTOz
4Yi/eXOzA73MoFq0dF7Bs0BXddH2YKHteb0EYKgBI6mv9BdAT+0PkpDf94VweOdnV4tHxvsOhlCf
mMB/rs2NLIKSRsjNh8MbeDyK/dolz/6Z2PAPQJMpCXTHl7ttKKde5csQWXVryMDLMrIoFtrHuvve
LN2Eek7Uwx7qsITxTB7ZLLIrIt4mcfQPaOoXQeph9ir5P0Gr2bzdXAX5nTT1Hlqk2g5v+oLPDPC0
0TnP86WDjyeUU7D4aFnvX9LRUtl7SgfIUJ1pb9EQ+MLpKIUTkdfq9RdDixhr2aF0py5I9UaKYPVg
ckSNzLBjSShl9ZCqd4S0ub21d/665IIsYJLweJl1h9jgCih1R5swm8rSG6R8M8ZRVBR3BFQXbm4c
NC3062SLNl5u5dV3PYYoILghRLA2by/lxynrsbDaJ3SXocUowPHQhbkDx5MkhewCjz7dQzXQDCGq
JmJohlqENzJ2D2Pel2/AXfdbplp7N2iWHhS74bmfncsviVTn/Qdz7RnZFRPzKoAlODwJSmlMnbLL
e//AFa1+9JfOUZkw7cHC7ZEx75oDjJAOwcYITWjjWa6U8I6+0wxpauu3gsM9U1MJ1BPE0YsglWWX
BMWGTgmDGhzTIl2aYPd9ymrFzOcNfGmV+neIbafBQlGOoCLlmcvObQLLMoeOewMUvP9YLdYEFScB
R0xCiVzYh4PTl7bi1rITtp97XjjckKgGVFotTRap8lT/arrax2/o6xbigQhv2E7esw/961RHqX19
Z8rNqTmC8SUcQylzrOC8NVK636P1v41xJ3VV4e5yrIzOcc9SALALSdJIfv2VDRLrr6s72zuQ0SwG
ZkX06uLQYQ4EXCsID1DoqKt1ed4QIvIK66+I9XLwyPYHXB/6IFUP49vzwNPRS41G9ofBYlA3e3wy
YLoK648OH/PCQGYQsgYuj/C5SbunfOTD16vtMuAVRetV+URn44ihM0n6JgWoe9Z7dS25Y870Lq1O
pxojjR1lTSLzElcTBC+HmKJwR900Z9UYOz1GGz/46e1D5pytvtr77S+8UahOMdSNgwfw81P6aEZu
rTLKrTetjK0YlH7pFJlg/Jo8PiUA6Xj9Q/U5wjjhahaBpiaCpSuEQN8gXNik8C0B5mNAPsbaE2N2
05XJGvJNfitnfNf8pVWSARk1yfUBxWuPXiYa6jhmTgwXLn8hVW76+PgoK1zvuKQ462ybZuYb7xNy
Maefl8r0/l2sVaPoA/fYNKNrm/L8iTpTxH2nTADvha3pBMqGK1absZHuahGXUsqvd6XiOhQHR/QG
rxBdJ+rgNLeN8qkQKh1vajdZeWOG8lP+h/OBFn8MroTKHhCtd/5mx5h4Gsy3OI3r8UK99Rbrlo3+
wqqmcW2gl9Rwofhf7gHQ6eZb0j3aPpknkpxhTf0l5RTvbRhtAR347z5nGJzeeevzti/DtgI4DoOK
IhnXu9l4C7wrgCA2VlBUk4+vCKr+2gBmun2s3Qbbx0hwOK1j5N+ORXi5U4Os6AlYKxgdcL9+vucL
eeWSS3CkfxhlGXBhvv0q43YZL2jdjpWa+Rfj8Xzh1vGjUUx/7zmeera2EsUSkqv6LbLj9OfFOH5n
AzTSEOCFiwdomyjBrvo0iQAM8W3vPIYmavn0JixwsKvIZo1q2v+KiTF+Xnu70mEmgBgIAcj0+yYl
j+WxpgvgjEig9vMk7hSWVUZryaxFse19W9Y53Sx61XjTGEfbJLRWTNtyH4GLGddPeEPCRy2hfp2a
crm07ltrsX87SmMN3JFk+StQfvagxsOnvcxLHA3lPbgW2bxFjO/xkDmMdYZs0B78tkB886CX2MmN
cYs390gOpdYlU0JxtUeX7gKth6yTyiUBek96cJNkGBWaK8DTGxlU80+HbjM7O/KnkR2qbxbbcD3i
8F0D8+kC8ncUMycHsuSGH4A6nl9jh5zx3r6MX1mpzheYMPjWlLG20IDPXZqLGs1eeDZ+pVUtm05b
DxwCgTITg3DsalJZ0S5tTK3MDsSV6CQ5s8Gr8HYN0ID41cBDlk1a9JXQLodXtxUbEhvtWwr2AGc+
HOc21v1cy/1EtGr4A4etQfYu9uWfM5THjTIY3PsJgf/JYsxstm1R5OqqtQULJqIKLQEKz6ij2HQl
Rg1lvkyG2YQ752cRjqIelXRYU5pUSjNiBaEc39eVNLXZRgAO4QnVw/WB4vrWoT0vlzybptC8jKSr
rP3jHIFaGEpCb2nwldkv8MVSlE0wYmQssD7XKF4AzplOa6qa3/khGqdovhCQ58wlM22rXr+x4Yuo
qr6lwMEVa0ar20S8owK6g0Dt44sVDcMKzojaW9W0mhpelx7OFgj5+vtnYpqddlnMO8Ak1yT9NbN3
Zbr6uRoJ6uSUL4oeUQt/3CeXcz6ArlryWaB9zAHhNo9qjGv1M+A17FP+XlHpZa9SAvUJC0bs49KM
IrgpB2yJxV2pDcnhajnY2hAvXhZ575UVfUk6HtGzKoREXIABl4wwFalkulBJaVBwUwFwyOnSWLau
t+mtPl3J221/2eOuAxad0yzccR1wLbExHmtMLN3Y91h2xNxGVMbN+K5y8Eu4qX7KvSXmmPxakXdv
/beTSv5WflCZJ7VMSpUQSs5r4EBvwvg1Ebc+xghiplWV0x2caOy8M/am5lha5CVXEveFCpK26spw
09kzR/8D/k0Jy0lThQTOgWUumQ3t9xM/oibhG4LpyUKoQcsTeTLITIlLOP+hK35+DtmsIhYhr5GL
s1ZPbVPHYSPaxemfzEE0E9K3Kc7ru3q0m4K+AJxEIavW+/CGXdl2eptm0n60UPJ0xb+iKBBNFuAo
TlKM6xQkd6pbsjKzqZuELCNcprQ75tny8CUK9sr1dmwpU5UHxMswjo9nwSLBSTg3IoDTP2ugwQ04
VrYJJYI/VNLV1ZxSx2L6F0uq4ehU54za8n3LCKluv4rVNnJVciq/8WRQ4sAngTHR0rLFMA8guNdo
lcq+MogKzxSsI5/D9UWOXIaeIrZwn8Mk0V/BKXd24gONaG9hVFrAtW+v4ruPkzPNbsvPv0F0/HX2
UqWzEb9vUHsvN6H5Dcd7hQkGOztePODDSf+/DBt0X92+lMruOFk/8+Xv0OT2aYgYFrkkNDR50O6T
AuroEdxj12QcmXl2E3y/VGcQUGnIpg6XsCfGpclkMCj1izKxRbBVJub6bE2do6du7O3NN3pqCv/3
UzVOj8qNO0bi8xTewW/DJWtQz0r+AZ7Fpqkbj81Awb/DrPSihc50fgodVdB9GFe5tmLvY3p7pl8H
Td3nQNSIyH3dZcGgqbRgFji5FUglCsBVHUJGo8lPZCwevHxKXpLKez16PPtqirkan65N3ZkHDXGg
92+8aIWawyYe6fiKh0Utn6eCsE7gpYKZZka+pgb/QtPnMWHmb5sRYRFISsrI1OhN+Kpwm/d/4d9/
+e+90O03lPW02MA4OemA7Iv9O+rFo9AR/ht28pq8bGr+9SKALN2WwLXB4DmRmLcB1/4bGxHY0DFU
WbduygoF83Dh6FVBFLl3QXDbsS05KxV6VSvtdTHV2om97fItf2QF51T2/+0M/a86afrCBbfRu7Ta
gRFQWD+KTZo++PZm5AiPl1FEG5XtpfHSyEaA57vVvzO05C3AzSCc77xwQ0sw9wGbIz+77VdSpDD2
PChxDlIQ9RLfSejknMPmkfg1c0p0nAxQiyhxjTxctJLbxZ0qQMTNEp1FcmQXl5sQT69e394DY2B4
zthAIbtq9HYxw7Op4miz6RUTY8TpOQwPDDZiLc0bxO3m2FiN1C6Bv8OkfKcarchgBx3cWaLdu1m5
hjsIofAxMYUkdhJq8R5pO7HOgSgrzP0vxLN25ZDBGZ4DY8ptwtoYjA9d8Jk38ZlIwfJECqjV1Nh3
3RkNRScR2XFimrQl8EA4toVlkMpEHFd1nnJmnpujY7K6GDQBW7yj1IdyFsT0KwK4dg9umafQQOkn
zZQ8yPbKiF4T9gYET2sMQqk8In+5Mc1u2pwY/IxFFwn6AiLtrN9LmD1Lr9T+u2ZTMKm55l2CjhKM
PwTWwfT4LmU9+fS3AYPuLJ2OrKbsW52Nyb+08J4raiIlX7DQdF1LxKitNBpDH1/LCRjPWqxqWL08
R6cgpPnbacJg4Tn1FiV98UXZ0uVWkLVNcDueK1wQt4cRlOGpzPvNdhNqUtLGo5p4bC3vv8wpdVcU
D6K/a5J54HzRGWi/L3i06BxIa1BI8+x4Wv9p7b+qYaY04HWD5Zk8jbIw6kzkjIthhH6DnF9prnYm
b6IkqLlBwpYaJ5aEWx1IK8nVaYjq3lByIxp+kpOAkI0Ef8YJZ9ziJRX0hWkvi3IDb5WWCyqqNyh/
1o026qQiJ4qLr+9ZjDD9MKx2JkTj0L7l2tBji2YsAbAxHMaed1wYj9DUwLHkYyXqiRXTJcIaS4FL
TTkqAnc6HsQInEOBOqHkkx9vgseY1GDoOXSeem1UXM1ODIVgRxfwp0BRgyGnS5vMfPFHq3QML1DB
IHYb5avnTp/w1m3MoXlHhHRLyKz5wyYJcE9fmA+M/vR/CGIHws8GcbpndCBLHgbmPykgtO1k7tx5
yDQmAj9kyB6h2564F0U4j9OhJL4kNIsEj8wOX/sy6xQnI4hRlmqVeaP/5NVKSFx1bDgatl11qdsH
+dzlrgaezG8bXpzDCIlHV+XoLHqQl7KQUFe75SVaw88+iG7H2PI379KARwMcA30SXHvXMVLFvWXN
SALl4A1tX6KFHB8ZjWUflj/Z+115Nz+Po4bNohw5fOaiqFl95/R/VSqgRpBFhyXH5mOzc/zW04hI
L79a0RU4UC1iCca3XgoAmjgAsV74PMSBmyrO1cmWmU+Mw4jCFBd/iKpuScF/PTMjiGOy31WUy2ty
EWU+JUYkqH25WrbFdq83UT/vntiBYMpMgkHfEqPV+cDlBn91GavR2DVizKu6iSGNuVBDV3jgvGAA
FvCMrrZi3lK0cPpFc+mLlImoKjaMfk7e8oZtTbx8H2NbIDnN+YT/UqOK0tU/He1IfYtQJRT57vgC
PbJsCxXAk/6Ilw8XdYvfa5ApVZvqczWJb90TiWQGHEk1wO4oesamS3QymZ+CFps3nMI9gVGOlY28
W9Nbcp5QzH9HOLflx/F+ecj0g2K3t6Oj7C6c4BZIuXcsnkUXdLZgwkkuzLgSdmUhX0O8PnXg/x1N
qDJLzc1P9fUMSBYHrT8cZ2heZd8Xy3qbdkyx0TfCYKwgTKxaacc39o2m9lXwZGFtJWzhFCHSTVbb
+jWGxJhqjONEY+zQNM+F5dpHU/UPOfF4F3vKwF63N/3au5tfCrwqdQawoMORjsL/R3x+/3N/8aDW
+SGFa5wNjOnCWZ9yuwr814wg0HbZpTtpo5Awk77q8bEy16UIfd1lWtLcUjFmz0Tj3wOK/dscj21L
s1UfPrzXBEgmaBU6nkA3sKMOyrL4GHbQR1QgXwhD5Zo9eEZAK76/5tEbwI1BstcNoYke+WvFYO+D
XfbnGFvf1RZ4RjxIe5+Z6sEpFf0LftunyOjQ52BA8V3JaDiPb8vRPFPGqpn2CZnK3PlPF1KlFrOF
EvqpqCOIrzeFu6MvuErjb/D9wZYdWmoKxxgtAmGOO5IL6KFTu/SHmYlJf5MFM9s92THtwlwzTt+V
4MKf95nGZDddOhvLeFACVf7ZXFyV7g9zuIAXeTMaV9B5Aio0Jys3sSCup1PUyVOuLkx3560cizXt
eMXjSEp4J4Ju7OvmYBhyZ8+YXkHy0paZfQl78e0bW0nNOu61U2Gd4iR8fzky1GpyDqv9UDuUwu+3
gvjxdbp7gZ34+VCwGulvMYjlcvu6k+3lh+7ylEenjxSG9M/YP9qqLe7zaGLP4Dut1Zb814iCvM1K
e0msUcLQZaQzvLv9wE+PXJz4HeVjd+X27iXGYgMJnTBxcKr1T4HoHdHtJENK3DvSSa9m6rzfOzgL
WIQrKh/NdRHBixGvP84WuCG9tmm8X1XXhSzhF1D0VhCFr8bOhQZ237f7ceTKu5ICNba9E7eX5aWu
GUPfTeq/jdEZ75rh9SnChfG9GZn7yYEbo7OcWfEVekak0Jb+0XTTWFDPhzq0IBqEM0/wsfefncBj
0/X1NlWll440qOlwR9F7191TyA8GU+zBpAhBbPjw0bq5PfU2EhyDrZbvnabN2liC0r17u3PwnauG
oPgVgEixKr8ruy0NBBWfhILGxjR8Uz3Lz3XbX9l36HHdm7IlGdeJUbPQBxrXCiubM9W43I8d6+su
OtYqixay7zG/kRLnwsa7XxcFh8+u6JcMtkuPOhtCA+nkzON1qtmfduxkB/BSriDPLGmuWpL3yMZ1
lJBX4r/vPYUAbJiRLuWqagwRz3tJYLqBolxB2A3BWqHSUtg2yWiAbax6uB6ufnMnW98JJruN1cM0
8RfvAr94pMIoh5rM7eRAtyAyaZ6pK/36pqFLXXn4vyizyEoGGtp34aTYqSCY79oKg4EcwwS+PePe
FthCjs6d9YkHM+We+iavz9fyWMUXkvgclLO7eSdFadawVXfmxQLymOHnasRZ6nBZ8JtajKuyn4/O
u4eJzs9SLFmnJpogw+0knx3hlASB7+2oUIFjrwJ1one6uvDR6qlGv7noAS2pzvV/T5/lD6TcL8Nl
igEO0Nl+WRqlYS1+cxCP+hpXIUlOeTRdIxpY9UQ95P5e/6Khxz93lDwKK8qUCeVZY4SUFt28UwMY
IWlukT0EsRcYVfGgqCd7I3SqIOsUx3AaH/Z7zQUmKnc0B22FqH+qIXCKZTwIzDmH9oFz98B5Y0oo
IYn/kM4mJ8zOplZ4V7HBgM9833pveEMap+FX7YxwnD+C9ypWbG1YvKNItW3AeGXlm4eUEH9pLsVY
gSa9vagLlha/AiNcOWD46bAhTal9pwJpuMLyFtpLKJ5Ob5fIuDuk4hyimZRnG6aEbKOkQLvQB0i9
IlADp2+bnzBQOaAWmfvpOwv447h9k009j7Tws8/0Qr14udTGE0BjTjcFVOMoy2N9jWc3f1CtDHIR
l9ZrK9gNVoFFtUzXK9wiYC70u8mJV4g/zV0ophKWa+smZxQAnSkq/uCA9y1dKGN7MKkID662qnw8
o9eBTgi3+GHmqruL5JK4ueq731oufoR1mjw1t8gwY7h01GMGb/zzkc9yNZ5HlELaB/b45SfdjMBJ
1cOs+DqX9puohn3tqFIHSNCdpSa0mbmQqZIYCjJRF9zVc62qKEymvfMrmWaDjbR/7osTKxu99jlq
mEWuWUdg4QH2Wp3/lD2cH+nkOmlME9TLBcQhbhK1FQUC6irR6YisdBGJDUBbHZ99rFn9cLufCuCa
HIe6szWf8tZKr0aSn7DQRNVZXpdWPLfmoVVnduI3t1YU9e/+HFBpP2NUZwcIwndWZNAyV+jfvfc3
DoKb6H0D+Oe/47Btb16qAz1kNF83SlSXaoa6M6BQE3HnnTpbdupOx8hYx4yp17QGFo0iGnrQOaot
h3FW4OVFkT6FrncCO+cLR5UzTirD1ha0MLNyww56pLRJRPC9zlFkgIg6td2nU4XyBMKyRED61gKl
515uINm3HcZ0QJv3reuookrjvpJ2hxsfEwcmw4+Y1F8wzfmAq7b3+NPhNb01Bq788Dog1c+oM/aB
mUd/QsaJbvcLZumpvdd+ElYaMxWeVF1Y4b66F9fpP58ulvhjXg0T5KbD8ChoocDPr8YkNnAljJQz
l+CsVX1A8XixjHXQntGXAWaxyJi+eAfrnTXAtai0wxgr7J1gMZEAaAwfpijqdtbEMuVHpV658NrV
atsPGTbsmLCtGvnhw60tfydftqig3ro8MIuN6Hl4bNvGryCQRiwDJhhg0RpmDvKjqa1q7Nn+PyvW
etrId246w2nzUW0UW6WQEjY2CEGcckekTdPEmoIxLw55geOH1RvXUB2Fks3wgn9WIkcCTel0V40t
LWOITPY0qgwJyXOgm3QCpDisInwAP5QhiCrirANSePg9GVABVMR5ZKNJdtSRjEj+74YP9jR3XL3C
TcktolkgE6ORWWCU1Es8LAy+Om/9XZQB7lkVuZukjTa4KYwErMUQU8tgV6p/Hx3mH9VtUHMj6IXe
AQEC5P+oYLQpaWfpJ+iOLB8gizNIEGTL4qc/gvZhQ7Y3dnsdTvnKVIexkL+9micKddnrwQAwTQui
Q2dY3Ue9PrE8Pt7ef8Fdk0YT5Zl668usyLlyYyh49ArUigItHacJ4zT4MLH0IBLPRrJ9jq9/FS6o
mUaqKKuMpvhfW8MIIzQh9b/OvY+9mQpU5mW58kb/ifkvPsqvFFWEICM6az1LQJdxRfJdftsFsRs6
vQTrh4auhwi6bgDD1mgHbkOwGudoJevOeWAITDX7sLJ7+awCDdFZbEeByJbAQsnkB0DMz/BnSFJX
0S6rO3VstrN+y41dK9NOqeOiUalerUJy/bk34kB1sUIEMvPG+FhkcFV4vNzvVE1OoEwtML797R4s
aRmJJvueFBeHHM3dRFLk16Vus/hZ2Jqca0q4L0QYpcTbfoGA8naDk1PvnRDzFX00OrbO/ikbJS8R
bA3VlU7CAb8NARzIhnVNBdHTAF8/mQVi9IgV6XL065PzBjAV628DeiPGcvXyN257EytTJzqIiGTp
aLBMohdeB0HDk6aVkF0aZPQpdz2Lv39H1ir1Fcx2pnm2wUlwbcYgrSkQ9XFt2rIW+g8n0+SnJ4xB
B/6lfr0hx40xXysFdCmjO4mYTyOOJB4vjQqnLyXlPqqa38qlgXffIj+YKu0WU1fAkYdmIwiFHGF8
roQG0vvTy7zTB0Mx/a9Bh5FfhoeObcpnwjAbP0hy3WdZ4dB0kaGZ7QiZdL3anxhPtOenDi0kIbIj
b2CkoZ1LJ9vXLqtM2zWhcgq3ftbFrAdu6ytep1CSvPKFlYPmNQXfAypV+UmgPWvltGTdiytW/exi
SDdKfH4/biosPEIPIz3MppuD0rXT8geYfUicE00ZuBDimOv2RimCczFe+nSq+QBTN+Tg7sIpm2ym
39sN0BVee+exn5rlFWKHMzb7c4MPl4X9G1vjY/XWe5toaDcFlpy2N4cp/ezZk+CyLWudV+LNKTsa
ajCc5mAqpbP1iBjN00woaNucia/8A0/IKZJ2XqUUrsUnLVH/K72jfw++W+cKa+dihPgGW7cLvuAd
s3VGn5btbvS9mKL4OBp5WIC/MctQb6U3BM/jewUQx2oWL0EKqYM9QMP34U+TTQbYpviWe/B9mASB
HTm8eLlI7af32uDQW6yRV80Gm+Aa0sx6/YpM7pYzwFZZrU9h0z3Girlm45z4Mq5gghsXfrjeY0Be
rhueVciioXw4rq4eb19jo0AtJFbDwc8XsKpK4vPsKUJqAWTApMJz/tYNIu3ASx6IOQLdbF+uLOkG
KqvR1vJGtqboGwI/pmJzfPWUC6/xGPv4oVLcfRyp8Iilhrmqfg+7secNQEY21Z1LL0IYCTuXXBcF
4u6gMdP8IPhAEgcmfI4eHwPT0Or6vDlIZvdINk6qb2mvqr/GxO+U6w+6ongO1fcYOIxm33DWhWP7
wDiGpM9Yx/BIYTowKr9Q5wi+iQjWcpgFx5GrdHQTBlk9Jgak4UqIAE/tC/QJ3Dujm05LKeUJHG+R
efnD0vfDPgQnK2fRwBeLPyTxAkoIRcoovItfP7ZxMvslZd7o+36uYNQqADAYR79i5kpJrh/Qvolc
B2P9s7yPLRsuC9la2f5moEXjUlaOu1cWKAu9LQf/CX33P0HeskwzQBN/oLfg3qsRE0Sm8XAp6jvR
/iMDh6uEW59ZDhTmXpmr0N9F1r4lLppgJjcxMLxMmcctcaDFwxGbFCIPkpYkD1aJM3fmx8CDQug6
99kZSMHm55M1vIIsdC5SzxhOpXvL8LdfWJpZtwVWE8sV1Qoc3vFLscfeJE1skBzujeXufG6W6rpU
pkPWWtPdYrDdVhuZ3bnaY/5uWFgu+ufSBDVhAystMS/TcHrSZVdiId1lJrTcVKKjT17gKpc5Qd3D
PEGJNmUXnx6T7C8+GEVnLOJJGUXbnsV3R9mmOTB8MQmuwD3ATeM4K6VUbR4hA3HzSqKgh5iNrkTz
fKfmQrKGpFsCC6Axb+fH0LGjo4I52Wl5IcUZH22ED/VegoZ7rizsLuvtSFMa5kjzzeVrOAUOcT1w
4yYVCwnjK0Ju6Ed7mz5tHxkZngJaZSY1lRRHzk1RRYrAR5ktCeja4avSoYBYUferCCrfZ+xNcmHz
yCOKYZA3EXxZ3yTr6fVMKTAoEi3tOJunn9KhbG/FG4M0hlbPz3DRZkMf/lihlTg2JtbSn7qXGIYk
TXacC1FEMj3QqY1FpCSGho6+zF6viyfry01vE+DXQwHqkCJps04tjHbXGau1lEBU0MB3q2GBsWK/
saNlz+x0lPXbqBSmMBZC4tlbZEVanuh6tMRSJFINfrgSbyBJAPppM5ty7sChxwIKKSop7TrqQUoV
Cf1TEbqijHu3O/jAjA0nptuP3qrs6gNR5DZ48rZqXF04D9rdCvpvOYoxcXdsTZt4Vr5s3lPpcBis
G6XVCMlm4WaB/AmHI2O3IVOIAORAR5WPDDDGLlASPSX13AWTRUzzK5rT2n92k0Jn7zlhJorgaKfc
p9Zna8li7SJj9kISaMZef0musaXyMt3UMla01z0Ah2Uy182lxSfSH1BMnpVex2Kd0xLZCKGpRedc
yD8ymMB1jmQ2OXmjzdiU3UyxdZ+1PJfBo7ib5o9vd5hYGhJthyvcjnPqXtM2qpNwIoCoeOuVAXjc
n2qFI1R7eOaQz2IfNJtlo7aM32achiiviv2jctiQTPG3JUNxfew4Z93SdvlvGZ2a4zLDtQMTY7qh
hE2yCVBwLtOMfKn0fxN4AvA5tentwz25QCz7g67SYSZ+ncVb0NrV4d54RLm6HOZe7yb6aHMRgzge
ld8aRt0+V169rT6NMN4ONNwFm/XF47vLB7qsu7p9kqHz7jI/Eh9FYZU1o8EHmvM96PGibVeZF/i4
gjpiCf9uk5Zkru6/NK4oH7JAciFRdnM0Eqjdk1Nh1adOyLobhNtOwtqd8GeIsuMYHpm1RZ8ZbIM2
QxDYSycURsTaNjRbFau2EbP0XPR5lH8ggrIhDimFLlesnDVO3DB/W93iIUcXc8B+L1azsRpQWW+A
O/f2EnFLauWUAPhua6O12x/lqVeP2OGx6ubfqtmGpgLnwy9Mo1QTMNINF/o0p+Br6+mXoMi9ai7V
fuynKKzJIBx99F1WvUO4ooEaGEAP07jHFPUv9M4hE7cOPSbOB6NbKF0whZv+JGF/kx1XZUtz7wdq
RMMThm4/ahKjHhhyCJmQ3Xj9E+I71RVwzLYY8aHzwLBJqtcz3Fljjl+BRQuJRWE/e3IKuDgHwPnO
RQFgZlkpwhJwuZkqxCCeErwwK8Sstn0LVaDhhCXlx1TJhwMc4fOQx8dZ9bl5iXczYbn+t//JUdnk
k+LqXXT2BjqZ9xLqbjFX/5ETeDuZqyRl7S7X5le03HwJGM6mQ+HmmO5hXZNvctQfI4LdSqbgnROb
TkdMdtzH69EVxOVRtPKECCUVeVIcrR2+R+ZKF53Y00XPj1BRyT+WAk/+5BI0+pycvOjnGuWL2l9D
ZTIVpH2qI7D/+I9HCzLTO+zCP/OExqvi6zdaVQrSSIf2FFcu7TWO93JNkP8ppoFaeFVFnD8vGqoY
OTrbxoiQM9D5TBUAK0FY7HqBqqEaDoluLTz/LASnXisWCyeq2T/ztpYt6BTJ4dwy7XfDpclRQ+tW
LqdAd68vvXOqZdfLYgdtv/mT/XyTVR13igBGnVLPSW2nTdEukS4+wFBn1T39p1dWV/jzmgkoTjtM
bYkOl5NJRG1kTixCYJXEmKvvjHr/1k+opjHPRCD3IQb+5dEHvWCx9gPDvSoRwDtscU0ypTWxe2Ax
ukuz4/DOn1oQPd7znFCwbVt6H1kuQt6Ickq0nmMIQegce+hG+On5r5zS/G4kiihqTT3WcHyryUd0
aHXMY4i6fP6NaMN15pS7Zq7v9UkH5l0pfRMURiklgJv7N97MfKF1NngMIdd7jwqAIAHDgjsO8tX/
G/gdH7vqiPfc7zrxjCkFn/+78Hku9bh8KNnKxXO8qvOmTpIW7x9G+IQ8qhfJOpcItmxPwMuVYbJz
HVW6P/sWPmbzMJBLO6fdpAdEXXHdPStg219UP3OlbDjyJtAf+Br2pFoADoOKo5GVLEVonEx2KB9n
paYTIgO6F2CzBNaGkfZgBLcyo0j3WTqojySe/CEr9vmo2h1tQKNoemLKUHZVVHLLZHZuoKg2WBBr
d4N5SZzfncVcS8uLJbr8t858LEyKyYLtjF82LzBoGMWFlnWnz9ITqnjFqOlhXY7bdv1YtnId/hCt
TKXJmy+Q2hz1YBngetGe2QU5LFA0g/8he9ZfT/1Exc0UJqcKxbklQBb9JOgAbFloyXB65TPH7tT4
fzHK/uSNKtDRSAjQtFxTsnCZzfLDX4PFXrhTd9BCi6G+LUrw9f28ysJgHsTg8enJsoRUi1dlk96r
ZgiVNzkXCq78ReZk/XEJh66DVsze6eS4mymnaF8PESXbJ4dsAMRe1MaxpbHDK900j6OhMSrznA8G
MTqTw2gXr1dBGjNDvZpZCOGfqap6F8rFjtuRbiBYAseWmj7o/+Xn6auya0/AzLx24b0i5W0xc22J
KISNO1wj9Nccrn6Jsg4K3IZy46zdQm1T/SR/O1DHyrVkZFhrBTGrc5ZBA1kyf4ApRiHAvMgCivuG
pK3tbAliXiO58PQ4/1yuKHTQhlqa8Xa94HFyYgseTk0fQ+BWOfQNbDHpU/nsaeZJfDkeObxusrmN
Xsosk1R7pIEn64DYIoIVIoIdPVgGzcc00osYl7nb8SVWZKJVTOFPk5p4Xb8ZnLfh88+Gdcjud87y
5bxf1yznXlbTDM+hYYrTxLhLj5OVDL2Nl9j8xD61zqG4nRmrO1ldNDUBZ5QeINxU8Si3Z40iFjn/
DHGhzaSU2lu3UiXS/C+xBtAArbxI7QI0gP1KrB0J8tSinOIb71fTZBEE9IAoFGLXa+yE5foPSLka
WW6CI0QXpXqWOleQhRDU7YBcHbgpqZJ54yMgpySjtw1/NWPSSSURgk1HGluxS1l57GB45ZQBdB2I
iDrBy+y47/kOrxW8qdyyVFVX0/aYXYwRxrJZ37wylXeunR1uSI1Bb/AYNfvdK1+y6hN79zRovA0t
rWwJqsRs5QZ0g0nKFJivtgJRqFmqZMfUM1AYl3S8QOc1HrtJyvsB5GG3ceGY8oM8kNqpabA8fdq0
U1fVgms+B9/HBwAZBAfTFOvShokn6XX7Z+1AuAhRt1KcJaWM+cfW5ObtLA/8yNMF+KqxafXJJHu1
ys4dCTcVcP+XXx3cZvKYGlcyk+nfO4/irSw7DrXiRN5KowBTMi0T9Lxr6/imLX201z5F4/CZRkBM
Hsnx4p8OGQcWA4XQXyfWt8QVxw6E5BXQCp+WnXHXjbyd/p6MeNCcbhC46LNeKXE26xXnDptjJGEt
AnzR0zssMbB0nlH/V5sGudsem8Peb3PJRkhmmXoDbUiDgqNKLPp919iSQvTXYiPiSnIXLu9hgyuy
HmwFOUzdUv88pyA5r9i19nYBFuYW8Sx1aUKMFidliGMtywEBEnOvqj6OZbobaMkMwyaFswMnnlwg
V8DuLR9MMKx3IBOwlvWrw99gAD18SwD3FRc1ghV3jKpojcpDJ1+tG0mzGTvTdv/++jhmnJe/SevG
yE/NbgxdixUS76Cd64HDcVzmf1zGA7uyZm3zvG5uqf8uFzfpdkvteP1kfzloWIiITfUOI6s3UAKv
k5TSzo2fIPvWtjiDTWpRCkq2en+s+PqSiDcVvxRN72vknvRNE9F0eeibUhil39oZTxS7/800JfWk
Ls0Qi4px/64bf0e2hTPC72Dl8oK13dtNgv/i7ujfJI/xeNKG6n9bp81qIhhRwA1GjA8bX2za0XUl
mr52A+CSJ8aRQuMUDSxy0hdfH05Wofmy9QTAhYcXco3fb6gJBO7E2MNbQ4fgajFdvBiKKp8vxdbZ
rjfCBZrRDeRnSq81w52FEhURG3R6e+BaylbMfhs3pvyrQa1ZPSUy9ZxFPV3F3tyzTKuxRwe/2+A3
A97Pls5ILaUoc27DBLbkkTCDh8FqOg6BeEH6zUtNjIC11g1qW8qG5Z8VBQTw7wlJJVsRViz0dk+W
RWVrsM5aOQt0YrNUBieeU9vo7OXw4k74KPZ+BN55pqOdb4Kxda6PCYd6tLctOdc4YtSaB/Nl8K3y
xE09yGIWdcWDE8ETyM5kLxm3XSSKmO2XtY6T7Ge7z/sv1fuqFJbQA/48f6Rrt7c4HymxLyNj8UFd
A+KXU201B3VUF2vO2dKiHPYVVL6HObexgURKWUk7hDEsfDHy6h3SRnZw8u/7A1zWCtBiaw29ET2t
ixV02R6i7oegWtPEKEYefVv7Ss25xIyT4UkTUPyxThPiGoHT+xAL7fwF5OoRYTU5090h7zTG1osV
j1GtQU1J3F1GkNiqAEWBskGicAJPwz9o0Smxz2Z1FahFrf3ZAxaDHU1Y3q5GrPpOGRt/oT1AVCZ3
7xizWD/l48W3kSJtwWjrEewSKIyNFOTbqxjakaVrRht7mHWudZAT88RWRpLRWqV5ulFEwJyPBwnn
gRIsrEwPiUPPVJwXd8a8sOegYEg88Tt8Jal9EDPh6cov9lxbwxkOpR/0HI5SyGpmob4a+eGlS9fy
f7dBvGOLvopjHrg5sT46htz2QoRk8IZhXVpLAR9uYUcQ6lhZzAWDD11Y/4Alf4iK9dYh3FBuKwDa
ZDCRQ5LEf/a5VKBsnh9wSrH8Y4DNT4ea1zosYBYurwH4j4obPbx7t0jLLpWkXIdkywFXfz/VvZua
JN9DO36ouZ+kUoeHyYxN1gtLmp+fNhstO+m9ZQuccEXxyx6XJhJu3HdrZTViT4HuSGwQA5NXCXFY
rUEEFg4zijU8PmfFrsDRxPXnSfL56+z3k5Fpf9v8w9/4oGc/nATUZk1O/3RJyeNAzAxGnupww0Nh
5LAuDcXX/lraUeC6+TGqOlMphijdqWGYaScgz/NgagZmHy+hN+F66GmHlowf1IjgDKb2VWpST/rW
XSITaSjNWIosviLe5WptdSZCftoKpgcgQn1G9EpJERPKc55HBrcOjJR1cxA7iHWEiHSckeAejmFu
6gog3E2c3xtxXMiKb88fBTdxpbd11BLToGWHoVotzrqEynja+Fev40pfq/864+oMt6ueOiUpqJcZ
5qP7XOsxF7wo5Be7cDmpBFEzR0h0f/r3lK83QA5JxKsnCYT3kLp6AwoB965tdgPxoMX6UIdUwZOK
aja+0n0SU13GZZ5yuGruIz3FanK0IKEdMJdULzVlL4gpf1bLlve/tsgui16l+nzhgLOsCx430t+F
CXxDpsyaSy1AD6ykTd7Ox8Iv7xOWKStbrpxuDBOhvQpa9cv1eGz5XDDcnZIvb+vCMzfchZCPSfkZ
4NwqkHFQQSY6zhAHpYTZAD+3eb4ytZBiYc7eAJOZ2+qQlXQLlVmjLfr+70tSPl8irgMLP6G2f56Z
WrQR45c8LfuNbGAH1SYEN/xHg4OqmCWQNyR5OfYcjNmf1l06Exb8q41SRsC4zADsu3PxQZ3XEwyR
EjjIPAr7Vv7YBbxfYxpR0mIWqSvsOChau7MHAW+RSRkIzpzNicdd6dfEhR8UWh/8mLKgvL+KYt7y
1iaqSBzViGF5yHuXL66df1VbE+6fURrONxBBDIyv2OSjo6p/0csAhhHuqpZz0zvXyqhK+r36sT3U
RsTd7Wtkh+7/84EYYQv1QCqTZuuMhWgTGBMxrjQUbHMUCmD4MngVN5C/AqqKV0ccigwLFrM9g2PB
+c+lksKA0pC8FKPlvF2wuBsov7U1+RstSBNDqB8II0oowLzqr7H643NcrYUEo37aJYiHRVwHfue9
wmEoOB0RLUryzHxXuZu8pdsHbfuM0zd9DThuyAR8/G8Wm06aKHeZFRXs45Q74/h6uQefxsQ9JKuB
hVq2sdUWVOLtkkSk9TZTP3y7jy+QEYk+INDh/+xgmDFpOkKrYGEoTAbe2TiorDyAgdZuQ+ocvwcj
GazbKvEnfeq1LTSHH7mWszAOwC881QxN7juJz4YJTO/n1iMYcyfQxA7laW8zEMvRfEUdOcMIig8s
20O21j5CCP0sR8YTl/hIwg1wXPRCjNoS3oL6Vgg0fiCUAWsFTqC/2LaU0qhuZV+ntVqWU/ZNRc53
00kyxUjpdoeYxFj0z7ru65dYAJ/CHexw9FsuGM6iP1T2hArm96t4nDEfiLVASNvLZs24qbIyW6EG
Q9S1gwMGsl70wtnCQPqKT0fpVXsBgyMcffNZo7ikwUxlrcgZzpSPHGyc4zYBS/0LcvZ0yvdBqUza
1dx+KMD47cOk317TNenQc3nIcAzjwKORMJutAx0DrQlnazfPBT9yYGqOF8pZ5TF4Z8BPNGYz0Ibn
8yy78UhdLSWEa66or5U2JNMMTrcZxBiXzt2O8pwlrHIjaNp+xc/tLuSxeZ94fhVOOc9KPkU5YH9t
fQ30tF9BgEWSDYOGdmlHzDgaAx8rKVB8E+DuFVGtWrfdiA9P9e49wes3uQbjK0fxxsmHRMv3RQXe
bnHz357itojrxJM5zg5VwqA/sUXVsEmPp7xyKMUb4GuFuJBfBRuo6Tkp9ahAVqhtSTXs64Q/r1fL
cQwbabMcM2/ks35Xgag9NLJDCHoG6LIpG4/R5OlnND0x3NUvrwW11vLyIYbnYQAgYm3o7lfAAt7r
vU/WXO15jiQg2DpL4sADkwqP9PNLBvnJg3H0JBsa/eIrwKUr97GGSd3qS0O4HMtjnmOlgTyIWh3D
C1Kz0Xqr7b/gy23uyWO6dnShvfYMUMeCX/k3x+R0InyCu/tBl9+QZmu7KNEaf2SyPcrT6yF0gKJk
CLIEo7XBSnjfOt72XsJCpliUZ91KGJB9DL9jm6pjp7iKNqEPkRJPbT/ut5ZaoVY2GTF9MolAwYlD
lpPejnVQfFegfNTN9JRc8mR27B+7warZOEou6C/+FmZ4DNN7PgQaSEfhRGsvB4sT4S36Dm1aUqbS
8UAQ1CeqgLcJMNX6UpjYSnkFUgqgTXFUpzixqkZXI6WYVjPa805W9Rx7QId2VeBYcZCggVn6vRy1
PYGuWSh2KhK9hm143aJy9uPPAn3mZsUc28xlrWXnkN5Bg0c5dk2jnnYBo5gJziH5Wd4wBi7WqEj2
RsWTar+FhrbGWhrhfbEVRzx2quDCFSJfoX2DxRxPx4Dg/V2yhdv89vVR55UqbzMOSyG7FrSjwFFk
aEjHcRKi3n3UIizHBrhpI8Jp87+0RnqMhgUrlKQ3jw9ypZDOkq8RdsF1y0AIj4x69rXfsvSio6D3
uht9RjPxPsnWT0KbQ4amZAp0frdTga2x5mxk2OLxLyBJjL8wWHWkftiZtAPX8va3wk/fG0dnwRjt
Leyud4I8DQfNKzDdXQ7eOJpch+jBpAC6We6v/M8/DzxLAmqyASdQ0tCQyGb/nk4JGAuSD36FlF20
fqXVy6iDdeBKURlJUMw3ZvBQBsEMCtJOCRA0pVRTucTMr+n5qbq2esar35oVyVrTPEvOXVyWtQYT
7CSt/w7IHxr0+NwsVCAnfHsfhK0wkGwgqucP4xIuFEIMQCiyn4kDd/LSNJkLxXSAK1SgMilgCANA
qRNZe0vdlKZ0iH0dC4tE4YiAfIl3Jh7I6BjIcA/U4xnWMITcSau+IGqBzIVEQ7ZwLOuSHMdBFCuh
lju7E1aaaRaeRstVm/3zUjXDkAHUdM5NAUqZC5uXVYZImw6vAuL5IJYvBVEebH4d8fKYXqI/N/fZ
Gwzfqa+IZRGn3E3N1nqapDGrMNf70/pTmT/DZMuSy8Nlg+fo/9Mq/kkOY3rNFTU/k2wCaBiS1B8o
UN5fGOavcRLaB+guCt3q9f3UzC49dTuYSzPlbum0hAPCWuNKbn8WfZGtYZjbo5/4cnVAICyQvczE
43CvE7yXYHaHWb8SQo0uAUGFfPeePrkzx2amUfIBm8QpVnnpNHJM2g/MNAyd3VqgC5KfP68dLPV5
cIxWYCZhPM39NQiQjbYbnNvk7LYqMwpISD+n3v/fBSP+K+PP4cSPK0wKkmrMK/lL/IuXxwKJECGy
LIAQZKx2WK4eMFjvcv6gdnjHvZ8nS8O+2SrvoGO9lByBMjWzXC7+ybQhPuNWb+3LojnHyXjJGsIA
AB+ywoWTJW+pdGyKlynggwL5SakyoIVkfmxp3UM4eHdAubJyUvs7V2l23XG+U3eNbX0KKbOV6EGl
m22SNSa7PrMKyAq+smP0gav9dl5hi+GOe574rGLSvDVpE/Lq8X4QbrIbGpZTu+uYGyOb76Dxu/9l
AeswJmjIitrSeYYA/aUVsHPXbz/wkZX/NDNNk9MBbJ2REJrydLg6xPhhcP0ac8tgCjUnjuVBJVZL
vPzCwFRQbSY4jILpG97rEY8j9hpTvOONorzNfYzGHcjfm15hok3cJPDzY9nLlS2uI1gwTp+sMExS
MVnEH8VgxkN14BtAlyrRFgPK9NzOEm4rGDfNwYGW8wQ1z0wEsTSOBlL4xisvEC4Y/SC5hmFNtuIR
zS1sDG3/gIr+DfsHdT6eqblCJ1c2rnN3Q6tuGtOhy3gf0r74GB95ltiRWwna/JwD9FeNu5quHrxl
NS10DPLqIbdvRdat+V5/HHiWLNUQvodh3wFhc0Xz19WfxrQBzJpYzyqegG0vXRpExHVtXyuFX8xi
UpoAJt2s5zlwxUqq0y0CvMZuGTppOdzlhqBcrJkw+0tMTQoe4DsFpCuaeJ+QvfsXS5VHVgELAbrv
z1nd6uYMo3oSLQJaSIPRiY8yW1nvR5uvkvzrz4Tl6yk7CcGhrXZ4LWEMKd3/LfHHtVxxMXiZSvX+
IVYcEwL6p44KfC0yjwDjlBfFkybrq02jER4p/EcxDK1WCI9ex12dB9pgNy4BiBFKhPFHRrr79PBZ
AHk1qQlYXZIbMUeXpGF6N+XaMReJb3UB2BkX1f/srrKW4CEmyjPY364IYRiBtv5PKXp2JusUfQ7L
g+uAKXeGd4+AoxuIf/4WiOAw/DvC2Mt8PAySZ1LG+OMyxd0sj3b7m8heYKSGsRCyDZo+pSIbcn6T
qDLgtOSWhDYsNGuin42KjHfOFiufU21unHaoBF5XPnOlf3awhOh/nO7uVC52gcNJlOqKo2bAVYNx
twy1jMmhxpNuV71FSA+u+sTm0/GRHXNBLPnz4fCaumToWjNstEE/5Ud+aLjKAK4U9fTpL20dYf77
pneBpMJrqhW6e7/BViW244WWZHBAk9mqigLIjL1wWVUMAMAK/WHy9AUNCctp7hpuZN8ueI6P7nCP
2J4UFm2ZpyinzHBEn0HV7YkoZ3Ow9/Z1iIrMM6h7pncI3jBBEztzIXeN7doEIR00IuXhAPTn0G7Q
lxSQwQVI4pXZCB30KhnKlhUdcIpXwtJE6cXU9lbF+GyTIaeSv/B4J6oYuK2/UPtPSoKwLBJaJwk2
sZoyZSt/umAd7cIoI5/mgV88tHsC4+1IRzIl48RqZKC/LsON1MZvPWZL/Id/NVzFOULNAfgqpuj0
wZ956yf3d681COKNLQ581lyObXP3oGpNe6eL4RQEULvyLQyHQgsnQmUYmUKFoACdhjjPW+F3nmNn
+sXkjow59kmYKDVJQbYv81D9g8G5eYw0DT4i27EVUmFoUVdYh1SyeOw04dtcONuoaaD1NPklSGj+
CMpWs0kSzGJvaJ9FC5A0WLb1OvsJOSeo2T70GcLzB6UbrY90AS9Tyx1Inl/zcnhsLdb9KLW8ohi5
2R15qrGr7GhC667iXk1q9g7xB/wtEPOa/KpoAgVGjTb1jxyLeAWIxJLIOkClo+ndvJSQvUtx/Gk7
fA6rCvTSYNweXp1+eBw9PQrvTA3Ago7Pkhv9N79xCkFL9mCbIYU4eNAuFe7Gbg6vlpElk/Uv4X8o
mEH8JQcK0bTFRf9ZIH8mplfl1Gc/IRBbPXPumJR1bA+qstr2cXON8h7HQHf5y/8Jzf3p/R90u3Td
dxx52SK2+/6dnqVrrNo86tq0bA95vi7pR8F870XXureLbvpsHbrOaCTnE/yc0vAUAFBT7ZWUEl8z
4N8AED+oQNQZXXqPfpZg/4KxeHWy522mjjhRmLh/CQGo+8EA66rki/rNpmxSXGiKn/S+vUULVluh
Fqsfs83aHWJgR3OXkp1SwCPw4qatOcWnW0DBNolH9S1ipTK+CceBEwwnBTP4Q5RHZO7dEEQhlCKK
7ELBImfrRGAbkKqgS2ImWHPr1gqV1rpPdrzEKTWysN+evkx7oH/BT2AV1h46eQ7PK5nbQWPYF5P4
C0PhKcUhI0eKEm65Q3s/jWsFW2cKeT3fjuI1WaVXW4+5QhEqs0LPUE0BkvUVcTAzQZNaOzZRledk
wu6LENZYoy5ar8Ne9HmZtRuld6q2oYvxVwPaVgq1gZv2aWlB3dmcUhbtektuPj5NgFq1rWFJupla
YjfvZfRhkDEfRu5cuteRTpQ72oAXJdYphYTreU0IUkXxRQ176MD1jEoNCguFUBMAXh3Hc6b8kqAL
1D817GE4+IXR82M7KgAzCIiubvqjC2LY8qtLuSQPmd+DYXaZwD0uRT1uWWmaeOblfajgDMVTnA9N
C5BErzf5vd5MBPuJqM32KcauEzt56QQKKKYwSulz/S6YHdSBSJtzY2srTSZ5I5MMiWOkgAnpb1IF
FLgi5taiJ7mnQ0exXODiOKn6JKOJLvAnOCii3I5zLeZiQ/UBleuIKxoUgjyvkQjKxAltRUcQW+BO
kmme6dyh66qsNFe2VvHBB546YuDeFDNsd/267L37vmSgZEljDq4pQXOujj1rKhpRyu7QbmH6TAed
QwjS4vYUfJClLRTK9pGCFpsh4a1htR63bzScifvN8qRxgCUJTFqp5nStdQpfWI0Pn7fFVz7EN8sV
30iR7KjXqNRzyVSv3tzTf2UQSyw7VJai2YleeiDKZF9QV6dr1RClnO+1am78H+LZfLwTrNMWacOa
Omy5h097tf3NWnY0gQfoXXEi9GeF0Iz98dKRHOvVHFEgXnMd+It3aIaCGganK3Z4MaIFEvFhcCbd
u+GREWrR+dHZ9Etjt5zK2u0VmwFe75mKyKFaUtbirOfYy3FKz+E3B4U1tlXYlH15ccSIq2SobClt
wviyp+MgQCSOCbr27Nn29DMSIK8KJTdxdGvMRqIQZ4sJIXE0Hu+6UpsLObx9vABr7OiUHIQv+yMn
yc034kXmwRJOWdaNNciu8rXBr6W7BxFP+ky7rp0T0XHCP3C6HCdp7vwYZv+b01g3SdoJGXgaeiD4
nyX8eOQYTfi8o9elXgQjdl/dq1/+PHQVE7RU0HC43C9da23b8CSk9q6Txie5uLpCj1UgJ81kpKcC
VcRACYARxvQhTMT1fwxSdNh4tPUBUN29NsH1rbvYtM0JF3KOBNhHQCts+Bux6ssZ3ddxg/RXvJ4B
aKQokmdoVBLZkfJXzPMQDzM3UVNrHekt+uJczOXKN9WfXZHzH5xsBeH6yMZWK3lHUkNHA32wUpEQ
tVJNREP9+owoVBDe7QXCSaUk8MTB+ENpLXpnr+CNuXvQbvr5+B/iNcsYLY7yKCcHKmbUo2XqtnwY
nhuq0xaqlpmoQi3bfGWX4NQhEnYpi5YW/lkP4wnI3sWL8deO29clMbp/aSZV7fXjXngOPmyjlEpi
q4t9kN+8sX23PTHM9pr88xSfvvrV+XYM3KLfjn7x0IfXoSgJoADqBgF4cVUN4yJFOJ5YIpzNrG1D
XBOsGAIA6AZQhP2xGtLvQLVTC3uX+ZdzC0fCrDSIhGAZgCUqzTifwP6D/2jZ4KnDSXg+zaY/er0G
hptTDAivEyB1D3gY608Qh8MQeEcYLykQD23jiEN1nlcpbm1a57MDkC4Wq9MgTPlFm9O3D9h8Xp5X
X2BXMCTaayykOCKjsrDITezQLoqzFfj6hUVcvzR21or1C8gnmB3S839GmqtfCR/gJ0cEYBbgCsKx
3bYVajO9fJvrUEibawMyoKrn3oTSNSOHmlEyPdk9dkLTuPL4plae377OPqpooS8FGIOLOPTnY97C
BPrCSGVJNOPRpxTfkoI68/qzC1WaEypMtaXoxdHZTyNHoVctq6VjtTBlunCgSmeh6aIXgWZF37Ae
jEJVk0jV0ymPf8G/mldAuuiJpPU7VcSXic+wXmqdjWpL82N/0liSezqrR8BfVimUf3EfMGFInbNa
8i/IhukPXph7DpzqDFF+uhv6b/86YFjbqDjwPF1QqA1od8R0Jia9uWshb95MyGMtwZB1rHUVbo9M
dnlz2EnDGfLew2K/FyurVeXr5OD7m97WvdxzlgYlRV+keY7fJcEHd/Ua/K2MoibEa0KkU3arFAam
sxPziEakEIotiykzUnzAoPbRnqDneHoqrHSWQuhKW/KZVv3/noHBKSAUQi4/7agsd95kzXScgIUh
1qzm/DuJrjF95PNz09j1jOMIw3Yy85FgxaStTPwDz0IZeH3eV4OEsFIy1QfnDp3ZeTqJcqwlaLjC
gy1yUtO0EewSI8B4bUwjFuLORkIp4tVMVuSh3RsLIxn6B3T7FxhzkIA9K/I7xRRASkxUVWv0fhau
v64YZtPBEGdmfZ+TKwPLEyIsVnMyn159KoXew5vEFZR7K2l1SK4SaQRllrtasaDp8kayphQ61D2Y
L+PU/PzOq7o6rcZqXiIm/CHz4c0p3t/qXx6q1CnzcZ8Yi+1hz3wDMjpzRByLuk1S6g2XmQxU1LsO
94xGd1+oJGIwlT4bc7vVR+H3OWjZ47X/Ybu5HCbvfKSQHjgwtOPruaMSK4TFgeKv82X9BdJuRfyD
ys3J7ekIKCcOa8wgGWh5RF/pjvixe9h7EO5wXVD5pzlpWWjOl/jROtfn7xbU7NdvhOeJ71DsALMO
g/moD3kIebc/z9U/NLz3INSgrRoKBtn5oc95wnEE7yYSJouHyOFMH3AsBUP0H88PMID6pICD9NyY
/j1Q7KuB5VtMo239xWdPlGBupJpCVOUTl7Z5Z1HeEk6Hg0kj2++MPZvWjBqyHG+tJbVMwEf4ig6Y
K9aJ5gGE1b5Z9egh/IJMuC/JjApl+fa1kByzSVm3q98TCC5ltUYiJJlqWaFq1k4xh+vGCoc3INaF
O3Z9NO+AXVfFS5YnhHAKruD8TmnLdJsYIuFh+EdvpS+vzzG88OTyTq7wgpCK64tJg/L5ymcq5NU8
zAnYmEWK6Wwd2VGEVhTaJQhE7pNb9p4zlJd+QZaBWkGuSb1f585CWsF3/aXKsHtxjaOUddnFxDqM
jxzYg/QJkCpmlDg4XnlLd0VSMTOOzJsRYqQcdGRHSzLIco3GG/AaBlKfedsmKrqPrPCPfvzxaZ/D
UwJCI3FCGI5f1fkiGrv6U5kAHsr8S9VF2dNLdj3KKUZCpz8Rqyd+wpRAxoTl3Mpz0ceADGJ2JQx/
JVTNTBOgBlhpFvfGDAcWD6dJReUZQSP5hFbniHmzN9ha1IMjwEN7PQrQoqYyUR4iz8+sPYfhzGTI
+PvMbNP6w7EaoUu19dR59ek6b5qSt0XuzEPBE2UZ1vcIrTiC6bq0dYzUEEHSl5vllFYUW7lJHZnR
8oIodQNll2as1gjDMlc3KaJb2Hfwy0eM4PX1mrzeVqDYNjgGAEz5ylBbYJoA+RNSqCS+60mF/gkM
dH00bZy5ka2MY+BaPpUpBQwNr7bBozUlr4bCCe/PKbrwN/WOjn8zf6/ph12UGF5o1bvG+/NIPtl/
wWOugghmP6GLMRZykPvxMH5AyAN4DZNUcXdDDzLKc+5DkyZf4A0mbOBAo5nGRq/HEC8hZZF/geO+
P5U2whwdFHPbCC2NjE0FhQAHL92JTL1obxxAYB6P+47fpBz4bAebi728xYrr94h5Z4WEY/5NNGdk
gIweSkFjFxUSqwZpf3XGNEz3wataJa3c6LTgk+6iavzxXAp2PSGrrAppmQyMLGH+6TxcadcaOgYe
GSHS0GI0QR93asqM83vBXh5aN4j57Ga8UaAjVGUv4dmJk/BimqzYpJ50To6aCwfAFWUAfuFnmsGn
6J1QZo5HY8rIRK88T6C0YtzOAB4VVspiFEQBqC6GcEIXo/He5yLEEKhmhjx/h1kQG/tu3t5sktO/
c+zL7CiqqH4TBcxiGpJ9NtQjkCdodE6hLqyrTh/TjOdU5fGAeihx6ucMUeWWBMhp2FvxLEIsbVs/
BNjtIO2iY55q8DDc3S/plx+07ETfcIoQetdWwSS39yvXFuhRULrLl+nkZjgrC3eZIYtwgMZoS2A7
m281PbzJgql/AiF6aalNZ8dREtmYKRqTsjy6gSoVJDCvNRt9m/q+cl7S9vOz6/sChacsUr4CBODb
jQYLITYP6bL0u4/9l7Atj6dfDsOYzxWVqmRazdWObWFdEJM2azoJzydSgC9mi31fz2va4UqMaHC5
9yzurQKs5RFapJL6qmltmxPYsrnObA2bcc+hxuRbGixTkJZeUyROBD8/R0gwmXXQ3TH9ThES2/Vv
GP4YHEP+wpfQjrhIlFB5iPVFsEzrwWfQMWCRYh6cyF3s8T/g/J2v3fhxHW3f3FuInjjbKVXZUPud
sVHZwo3Gi3RoToFzvk8Kh34gcP8RiAUGEpTCr0ikowHh27L/Pp4OU43V5zHoFhBnGyBdnRVgowvK
CDQM+mEbJwqNC3vyYinFnCEhCSLjQPoVXNss2tji2z8bt8IkKiTbeL4EU5RmAuFEOLGl52efUETj
1LG2lM1ZCtpgNZtzTb6tvWDUrDznSyubwlhe6kSMLhlQw7hiv2lr3n8oT3HiyDi0jO0XsR41K1dC
WOGm9anP4M92AaZqvwwDaYzG4u6psAz4nhOj/nrIHZFLlkdf6T0ltntDc1iIj7E7OVl/InMnQH0N
7BpDVRVU+NJZW1A1V+uzEo8uxtK0SiQ8kmM98cceWcP881kn6Eq4Wn5sX1j9hLZQzZfvoR4krjAM
0RJoTbhAJh1MFcMGOPOwSKsPWJHAOGMRXTvAq0oRKSPDGRuBbPgviFsHlGHR28ql5mUu3bR/2IB9
uyygyxnpAq4XRypjAKVUMt6LBghjppKIP1f0uVJhf3KGDaxvtH7bKbyoEk9fl4LtIUoao6pOjj/y
g5WoRyKCI7XACCk5v3OLWd49IPch3Yt9u4oCZ+8JgTL0igd1ygY1oagXoFkO7TptY904akCbYTOG
Wk6+9PZ6uP47WbvN5jkyKkQhN4kMMgcoKaa+bszFi+epfMz5TJIBlT+di+GTwYDItB+cGTmK1OY7
P1nTxePy6iWThFDc9tcwfUdgD5ae/3ygFwjklS69/dQa0O8VaTsMk9pegQjXeD3bfl//M+Zdfi0b
K7WCcfjqh42w8ytZxs9X8mUlY1aZtaF2igE4H8y7mk0SmhEIIxM5ETeRH11MtUY9z+n4azgxm/l1
hQbEnNyDwSc9qCkZqeTIr6Dm/TWi3WS+UVMinXkLqCLhlHFbXQBXMj4NrTyxgQ/zfikn3RJGSSyb
BtKOH9ts+F7s3+fRmu8uGll/wVCDISiKIaA/wivylMpNfhwnL1LBlqBIo3HcrGpC5KQ8yB5N4XCx
I/P9Q+/2bF5H4iD+xbnWE5eZKpUW2XWB2B0W3Sa6vfCss/CnV37ZtJE8guXv+eHhowbjFl149C/c
UaoU8EzyqntpaaZdtOj6E+11OW/wn/Xb77UMIL89bHIS4GszeUfNz/ifKkhJj0j7/eKtb2fD+Fxo
eHGAwPeyOH9I6RVDhnxKWBZs4uM0o/aBTl2P3cRhqJtVp0a3DNTwYKRZRrrCiAcR3PSmK8sIVQbS
3hHCk4snEw2X8reYNIsVYjbPKZUNOM+QG5wJEMJQq5jtc/BpnajXchDiYUA3QBkq102e01cnAj0E
wGYdZ8ZErnGD/BE6mfoTO8T0VxQXziHmXsSA0ToLDnmRaPRkMMe8efJkj0r+EosuFSQNgaO5LIX7
26TiUF0R6wnEIb0MGpw83KcYzKghbqMMfYoVT6OOazZLwm6g7ASG6cJOTjNkAH2QtbwvidGywbMN
9xn9SFFCXu9xD8H6n2YvvhUOm6PTrk//01JeVYYuVQePoU1i0NZJnM/1uw8ASZcyvpx3vm65aq1r
fSmUOKk5/6jQK9lqLp6K9z51bA9dgOL3MS1EdZq1LBbfCf7zRixHm0BLux5ST4WXRwsTNaEbe7Pu
iFk74koXGEJDix9Cm3VdTcTu64CzYtqe5GrPXCatSY6XO1T2ZmSabTPvXMjaqylQvTOoWw3WOMC7
y/C9glbNVM8vuW4FoQ0uNnzVWl104Jr9sdlNgkEwTLVLHxqSN+S1FyEFa8NiItDs7j/Gb20WH+UE
091/bzQ/gF83yYCmDJcUaJxxFuAkFXU4SUj+dmRao8jPQI0GgidViYCf6tDmJ7ZaOBK0oadyzHtr
Dw+A0fhZim0pCJymRxk1lfSxPPecDWU/5gJmbfFb5Twjf8jEWXxKOplhsTlj9uNmWHDBaEeIBjIX
wl2PNJ3yohg8MvvIrWzpVTo4YCdlNTOwDdjKP6GNSqZSL1r2kCrJP9MZyQkPMMOUIeuelMWTXYVn
dJSQ7Hpj8azsM4VQtE2GnWZIoUeUSaXzY8sXDUUYN9reBUWqHGq79Jsp0MeB3PSIRJvCjHsEUReF
Xbe8tyH7lNiw7iU38NMcijPLnZ7aT/s5TbBnw7nGhw6CyNizyT0cuzzRbRCiHN5v3XIbnSscFdE2
DmMTVQ8KEPa1pgLHzN0M/HD8i3XW6gfFUxUCO6NAsf3QjqTsK3rqVBOqkKUmXoAjwuMGIQ138RlP
Ql/XX6vyGK12oeE+Xckk5iZGJktron5yIskKcTArH4utDqbtzGylWQDiDUYEE8EmOXhs7/Hcacgy
PkxHKiMCzzwWbotH6Y3LjtEE40duQTYr017WH17yGdgfFym5cXT6nhQhchWkMfvPbPAFEDz7TmFi
ryF3dP4YGmvbI98rvQpVmOpTmqbt8jCsxsLkKe7wa6HQ3gn4L9wF75Ry5fGhN7YGpLDSOEKSCByL
jIKi3PbB8Sg7kSiN7F98euhnwI6af1dyTaG2SaSnGI5IswDTm07KY2wY+3KusBmyweOhY+ZQjHgI
mTN7QRe81CpQyT0cb/6Dl6NavsDzRSURYJOGQV4SsjXf7Lq5T0KxOaTbSCJU9CHi91snpYYE/Z2d
928DLkBnS01fZCUGpfNjNS/cQMIBuw+zjKCjgl2UDVvDtNZiSBDVbKbmrEzVAzwOIjxt0xkWhlLN
BrpG5EwnQu7Yk5ZTo//5I2Jymwr3hv4Y8rkhxEhbq8A1NhKmN7J0tISqzF8F0+LTXwZUN6nYSSx/
kPIIEtPzwP0oYfiQQ3JHATCItmQZkGcukCTmM0LEDi7VJxULSZtWWPRXdIAR0hkSDlh5IKpr9J60
4TXvbDzFZJbiVZoImxA78YG4G5b4Qk4P4wTF/jwdmnOtq4NErgtYgJDPyBMlTgnIHwUMdfx4a4Gw
SaHZwKBlUMXOoMTsbGyzk/KU7946UGAynwY9qyG/zaW7mhLkKn0G5GYLiCwWzt7AeISK6zmrTfiF
5fWYv9wgwRO69Te7ZnQu1CnTbbOcj/7ItAkfeenAvxKEPNs+cOBciCgkbrkU9DocIY5EqBUQlPvt
vB+no+iuCnxeLKT1Mq2I+4u84Zn3S6DL+uGSX9vCNgFHe/uweuiw2mWNGrlFdrESSfSPMKrXEoMz
1sPj5JfoeHEUkVz8FbSyNdxzEQabHGyHRfvrOKp+tKk5jMmdQmTVUaakYZ9mDMlf1qWzMeixpXab
RohONXi4aqcxIqPFZCJqCDrExyDWCbsbpt+Qp6HXbW80I97cebUDS1aTIsQsO/6VofNRqrGCDHd4
GsFluXJ34ZFkIsqlLjfaVx1JB5dJdbtWGWrEeEELXaWbOYsKUKFxm4NzHO+s8UU9odfmsXyPr5w8
TV3EResgKjil9tp1Y/3BgXoHxQ5nL/a5v/+kCDjir7sPHaMy5AaSpgY7srN0ZbfrTJw5yTXJ8LPJ
rgryg9mQr3ikYXCXBm7Q2OMSubJyufX+yHP78FG2BJVDWV5ZwBdgU3rCsmc9is31vfgBT9JYCBvP
x7iRXe3UFw3N+P6R8UvKdJhldfZCv9MKrNAfg4HXSKUq+YijmFu5WLCUqwwrf1P1/+FIbfTHLmGr
eoGbIxuo7ow5Mcm+GnMu8N8dgIUhueFN+gSYJI7VNBUE8MmhdPCcXDaoyUZbK4NQCXRND+cJzT9z
339g8UZhvbDNYTDkIn92vbAQaxE2qrt5WpX6cOn6llXxKT417wKpnnViKZXGm+gFVD3tMQjrB5Jx
35PjRyrsUKe0iJ3nJeZo33gImThCASb7HfM9ZQOwS2YBRZ4fGwSQZCJ97EgPnwpaxYwf2WCHNLUb
DYNiR5SB7rrN1gPEcdJZUxrCYYCheYDX+4bMWJHXHbGlNAWAgG7ZzP2m3ry2kAGtB3wMCbEq/PRs
x/4o5OlLuvmA/ztcxlvio6i+ZwzaB0Uj6gOPh+D2Tz50c70tyWYootLmmPtgZqzCcOE/NT0TiWry
+FQXaTw8brwxvG6oUuY2uvg2ir1p2VYvzpdfH5A2Z/CS1taeLbpyhaiCVrjJdXBs8Pl4cW4juRkX
MHS3E6chY8rpPq58bmtPwQKFPBLKW6if6S3TEvJRFn9/pIjjvsueBb7DBq9NtATX07qAfqnbrHTc
M81pL+yuDP4WCaQNxSVjNGZU9RA0u9zPy+EXxk+bIQsxNKFBCY3K5BjcAWeC41/eVz9jvfD7ptli
064sI0qDRrt7osCCigcgWo8gUGtfEbf7joFISt+wD98CtouKomMaLH4l74x7iyDajgRJ8ZcdtLb/
FU0NrIs5kwvJ37LGhoBIPRdcqAdYK+ymFurkw62uycPc8ORQs4i9gn6dpWkC7eZZ25Yfz/uHUuHc
k8zFGOM8ZS53MqHQUCvTIardU2Oi3dH0Vkbs5XftjKGQB4ZqTcqsKg1G4jf3XJ50V2nWoDtIdPIO
tdA5LlKC7KyAp/hlwhIkuzrJOT4iLp7aNNioYuW+IHwyR/ZiE06n0oK2dWeDpBWUHmq2Ze9uy/4b
PqgKypwykhKat7f3JjSyX4cDo1vzpOUYc244BhmZ+0gnSUmJt77ACj0w7j7EpYbG7hgFpnRJABKl
8jh/cRSc9l6B+WduWPPLACZAYF5+LzyzpBCaPHJl1ETMajsI8/HxQWrdkThoJwLMpJuadM/DpyYo
Tha71w/qeX7uouAw6PPvwIBnsHZV687JtK18GYBokkhsh20hs8XDH49OOXXGW6gCfkt5ybWkPSGD
OcCLt3B0Ssbk3TKiRRamKGkrjtLccA0p4TIHNQLQvnuGftqRJ6qxc920UyfUr0Rcbbjh4oq/Kalc
bb79ejcC0CUsNZWgTwtQN3aTUHlsTwqcoTz+mOjafFD2Rf82SKemW/ZZbPu9WumVaeLkOgxfOLnF
Dy6LjUA+ksFPz0i/FJMTNwYRjWq+qlHULo+fzE9zvN1dBTO0EYhHERSh6237MKybJC7kOzUZAukD
nhCNEoP2tMMCEjRJbPuC3pteD3mz1DRWb0EpIlKubxHS17CGFCsn+6p1fmDpfC5sBQ5QmV1ngWxX
nDM/AJZINUidPfCH7sD/G8y5AW2hn6wHueckPV2iZeZGwj59XiPlzZCjngJLN57FjJhlKiBdWHA0
v39zkhhDs0pdFeXXMcF1qFwb74hCbCPOpgJm/T13GDTm40w7PNu9SUy69lcAH3/Lp3KIQAaz1J4Q
3cWFVhuZYDHiJ0gYl8ZvcbAIsrDmwaCv21o7SRXnqzxdyS3sl6eVGa5LLd+TJ93PvHwfEqLHMN64
FD3O5glVY2pqAamPx6fLrehh3AeKRcVkFz01yzSn/Tr1TQSshV39bNYBEl6Dcw5gO5S7byhh3lJg
9ywpWR9UewVE+lKzwmqxELA4K2HNn6nIARHIi1idAh/pKV59lRP0+XyFfpFQ4CXQ9+janQ6/NsM/
xhCxrhjLutejijCPqXa+MxzFIkMoSMvBy2BXD9LzMSdKxu6T5jJwzJ0Jg8BQvxv1qrZ73qLr7GQI
PHSEhsRYMymvJa26ysvCA0z8EgkjG3kT0FxvNSlLrkrocJQ6pRotBhjakaW91P9il4UOZBryZKH6
7oFXXAo7XGKAFecSXiLcZcfSGrTiUFTE+uHJJ+n9AELiborhmmazZzOfkoZ9DLNmCLLNLvHSyWDF
RAJG9O1qOJLh+zULNz/TFp6GAC6Bn2uuIwGfm61Q+jJZ/VGkDoc6Cd8mAaIvEUVSy/MBtMU0ktCW
7uJ6Kha94ZTDbuPIm3VZSUaV5TwCDn9yyDURwLGkOE4OsQY0Kz+gKPFcDW4KNeovO39+CJ8GgM8e
1oqK/Adw2l8v9rO9UfluNZRM4+OLvgAXCdV7zPK2oTnPBWNKpZncc8W//CVLXaai2+VIck9QKH6F
MJVN645KCL8Jk+F+RNEs2uQZeb9RxYFtTRsuxaxh1PxaVinkoEFmjRwCx887/FgJ3AGkWjRnqzuN
RSWHt7LTlCFiBWng37V6GIK1B3J9kr4SxsnIP6MkaAOZPSoL63wJODXXpCK50SSl4VnkE4Lypwxl
jn9CEOnqWwgmiZ08gsmhGNC6MjSfb/VM37DVyMo8f1HYG5l1w705GeIGLUQag86+w6vzBbR4dBzL
VHbLMVR4iFDJRtKxU5r2RcL3v3T7/tpATWpWnbeweHo86n8b7xllrSyFPYaeoqZ6hYaYPZMYlY0E
50zWDeSRyrBCWIzXSxZgcn1Fd2L3qp/O8NcDWlYnnpTDA82MzIZANNQ7bvmUqwJSXAyLCpow5fiA
A0XsLg/wIjZI03Cr5gzhlRyU4D+nQYkkdOWJNGa/xXggy/9ILSYEkT56zoYHyTDIlo69SzP7qH3Q
Y3A2TpyUKmdR9suRfrwLhyCMqmv0gewzRL/dvSeO1eNEv67kyC5OUCMHLYgDKkZEKFpuM8Y6iuGK
+UntRQ91IY2kkZZ74MO2QQ5ZspiAIBfRSL1pVV/oaL9xxA+CtLvPZMpLk6bcDdIcWRBJMyXWsR1N
C4wmZ/XU/NGkIvbSFO8FLUjcUK/IdRz5CwvDKvME+LA16bT3c/0zPMxCnjhjA8cDIZUKrqJBNtc0
YCf0rtg/w8QI8QAeLRiC05Uqp+P3dH3VlF2ZsOCRvLHkGXTp9pKjSP2p/5Lbr4aTD09y2KOZyC7o
WV2h6ZJgZzVffA7k1A6Ut9UOuZ41GXBkNxJHDUPxgWflu7FjLXPNzNfbZBnxD6o2nd8fO+oUIB3J
ldEmgj4OloILwC3G1ihhMpK7TTWdWXwPNip4TJfEx/9z3XTNDTAR9LwWc/Gn/f5oxa/q8Prhig2L
FNhziHnX9ED1Hzqc/1CpFeuuMzfpoxGO9R/MKLPIJrjNLxQexH1ZI4p+B8t3DKQ08om9nrd91h8q
QWIz+69wZqA9IHv2x+NB/mS4wwCb6ILQR4yGUYIQCs8IlTm5YkNU+WSK71q2DNQIEmWZq/9wFCef
0NNLjm4e4FegFmBTe7zPjl2CZo7QoO4DnViwojxPUF5KHF0p1xa8ieOYkYM/TDxuY+DefrQG7N3+
3jeiPcNgYXF677A5YZ4Ibk+bGVDk/JbU+gcGCL6r0dbzqHTHONxMXLJUV9+e8qsKnHB6tdR/Zu4Y
BxCVhEVHoQCg4DbVKrj/ldWPUtfsF7AN7w1/7HuLFDIREkkDMLVtEmwusbwXAg4FcINk/9T/6plw
aAfaH0OHyYg/UFshhRD3QhSzZ0wtiacaf45DUUWrMXs9gGha2JOPxgq31qzxi8ttHKY5B776Ciun
DmVAi9XUn8Ed9TwS2LUcsVXSskaVOyaKmo8KbrCxIfPW61DhLE8gOkUdgF0tTkkDv/IpbjbffMM8
+fLFEhmbTqnrno1s6vLLyuCPD1UfBKdZOjnIYc8f+ENhl+BKjbohRcCMx/SY2PHiXjhrGoJrTNeo
M1BayTuaFa5RCXW4atAerSeKtLtd4GzsqFOCNno0jyQfFk6og5RPRWty1zWVPTjLsx6Yg/Dq9FlO
CbcxPxFJ47ey29EZkyQssism5rvt29UIS4cGHGu5mwNY9mtrxGCGrYmwMEQXoMM3ZUzZNGqYQkeu
qRkUF0zBQPeyL2J/BJzutfYVs+FsirDyWdpNky11Gg4Y4d0PSKUrEQMzrhJLy6jzhIrlxQU6cKGf
rk1IrvJwi1E87JCDL8Le2sgaVWbLat+aE8Ae7/+RrVzORl1/iFGybVNNo5KkDEE+8nbq5+lPI2Jj
w8yJJQMX9CdTvmGjKh++g/UL/DGg/ZaTJorhj4SmvsPXdJ8fWttHHXrP4wsAkUWDuSjWDEFOxz7B
DSpCPSGoj56aPnqJECMyO3qyrtIhkmhLea4zR89LB0DK6lOpxhMcvmoFNhgiYVmED9r/fDoOZNIU
reCuevdu1GO1MBCjN5FjsHrkocyaGHPuN2h3ipv4ws9wWpR2mDW7qyU0H2YOFhjMo8CnDQY9tEke
VpeZ0FxxBJkEq1pvyGUHDQKuex7tpVao7j7BSEK5HI8YnFZCVpKvHZZfGCj1zDVhhvUFno/bAlUb
v8iYL3dLVKnixmLhJVGeWcgk9RF7g4MWJSGDLzgkE5bpnKUZHVHHG4nhjHouxUMnZ1QzPWeUMiLo
DfxH7JZkHb8haLP5QknGVAS23Y+XPWyZ5uyQ3p8g7h1uCtcTNQ8DzSUWNrZ82EUBuxxFo0PsvRkJ
f8dXKMKhQuQMdknob+OsDJ52oNwk0Og5OMbKZB0oped8JwOdKK+9CCQR9zXljYmsDFHpfWlZ7DuF
UHKdMHc0xKCoUjGTXBM/uzu1BHJ5thiqqrajawTKwOEFqESScL1w9iugoZaC20vWJb4LcZcRI8ac
uhDjaR6+lF+QnYM6V1jwXBCBhzk6FYdyreH4mdv/XlpK2hbadRKuIE04A8R1NuQMlsXSvhMf+ECF
0DZexZfdsV6j8ermumM1aDvC2+dZWI/Ko2iIYOHLG3xbtBXTGtRtcdqP2QgBZXLCq1IPWFdBWZSw
zH3rIH2VWWsTLmWC4APZ8hzMDtuapJFPdLGi2HUfbsshZ+O+rNNslWcRAjmNXYkOyFB1mQs4J0fu
lzRopeCP06uLcZ6GVcAJ3s8rf/1eeuDM8WPdLiqG4BeGzhGjeHeFNXOdk6hs7cl/F8FVqTv7Ito8
v1FAR9LoG/FOPXkxw1QF0e9BDtC4HsZjxm81Y5mvqBBch897HE8U/Vwr02nCjYaN2BJU2ooi/EEE
3oFrxyqwx0Gjm2fXgRma5+p0R30tqANqn0nhohH0zQlu3Rif9ioKS7w0ndsa4GzdYHZ7F0QMZgRb
WwAZqtfLooQnbha2w6CAO2xyaYk0VKk1ry01tPS70GvQqmCBja0yUkgsPy6hmKh5RypCqAeHatqJ
R+uHeUSWLX5UeqzHrrN7rc2LWlP9wuhuaBu9dgckCTahOHeBivymx/3nHbvggWK8o372z7W3uuNx
tPGMD6vheEDohNKhr7ZZWHbk2wgLkBA9dIoW+SuqfhYCJCtz5Ey1dhQkhsotGAhpCVKymwF645BW
Pb6bsuHU1lterLgSz6gBADalYSd13Seltetf3dn2qRZHh50yCb5oEkDATByKyan5Bp75Ypcjqr19
rozuPxiiCK2WJnJaWcEKOWFVx2Os0UN7gwc6VVSNZJ4AKZqtSP6J58LIl0ScfO9dKLZQC05IxaEx
mRckI+qxdsNUJPTnIEhnykOJJjWRqb9qP+VQUaZCAHMbRPsnUR4vo5Ah7Zjfy0F9U2zdR7Eequ/q
Q21RwKysHqz/smXXxkpXu9nqNPLApTGg4yuR6XC641VJc8e4KUGzYTqQVyvkn5Y02p0cJHSAC+iC
vjZP473kW2a/EfJv8W1NKtzz/YnC6ouzBDbuiCuHdllCN5OVPjjdqMpGqqMoURRZE5jXfgALNYEX
YevcKqT6ddi69VtP0RaqcYngvQLKfxVQUTwJ8kpjoBl9j8IL7eUMNawRTtdqW1mlU/Ow0v0eXSAi
6+v4X2DGKgIB4D2QRT2hCWW/j4M1Rox7Go8SqPZPqrKjOcUEMe5YXGSmdnN/5Pzxt97SWVZG93Dm
GLMBJUqltcAM/WHWT7wjUyjET00IFxnEBkS0sThgGFHLmmR0NWlm4MjkdiVQxCqv2YnjCVGv9wW0
HKixtmU4mHatEIobq7SBWg1ZkOg2l1uvmbujaDXRMr/yL/tysztE3HKEx8UAPKndZvP+xVsSA504
NsfsJ4WYy5rRKVtvrfz21pft+j964mMEaCxgWQ/QXNtPEx3V/yFlR0jZICRjn8mVgQIoeciv0NoA
y5Mkye4WLYTCUxMC33D4TyjKkg9WK2lGJZDY5X0FJ8xeM+sfcy5TMA6lLVN9RUKLFkguAjSjOPcx
gjBLyNTfa2wc0nRNXwiCF32/l1548xhlrO1M4ab94UMYZ+lXVUT5Lh3VFiEyfUZBjqFh8Vv8LSv+
Jx/guRtXmFNb+9XBb6d4yKulQln3IXpOzoIRy8rQdVk8brtp8x30nB/+S0pQ/3hqsjt+GNZw2H1J
XOZFyrFRuDQ3rB02gkeWAWI0uJYlOfLFCTsGKpTHRJ57i0B6loeLYqxHYoECfWpJUYGDpOU6xFYP
Qp0lw3kkquSEpd0+HFvpgz2rlK9MZpepSYuSxy+e6jk8AeR5lGR40EmcDUg/lxZJgY/i4CmjPTyU
wmLBs7uEahdUMzb/QEv+y16XkRFDMRaBgmgckOmZwiSq3uluwRDNZ7KNS+KWMvamr/cMlfOdSxkv
OApp9S+426BUEl9EPwlRS7FFqD+nbr+xtysjAnlmMFip5U43IbFfMjsevfTywsBnxc3ArebWvoon
d57SuI4PC3CYNDhNNDp7KWq5x0Y4Ge0TVnCncuwPOBWzIZO+X1eyotOMrFw+opWOGY4hPgLP5OEi
GV7Tr7290BlEiAH1cYTfQmGnL0QBDZsjOeigNcq+fPA74BcSrsdeKg5NfakwBCuQx77fNVmzl/Wl
VBXzH/3dgpMJBqdNKNQmzK9xX5s4JvcMdwkVhKMyUq+Vbw/dhX1ODHkCtnVsznEgznEHlemRi7GY
GGmWRmx6GqqIlrq3muLoMP02An2KWHrZSAmG6IhgAHAuFRBNtrH8ZVwUjukjcuu0NhP5/rc6LB1M
c/n0TODyvCkSClswldhwTKuw+wx+bsSJ71qpp2A7qa3VfbxcY9FgyA17Au/f309T3ol5S26Kw0+1
HkmTrH2IHiY4ia41vWCMz3ZpiuIkjBqcHI06q8OiUUNHBKTRuUoVpKPSMzltT9DjIpjRWMTIJ2HC
JrhEagjOyU5NqSe6K7yAUP0Nwu0DNUMMRctcC/8K2RN4BUCb2A/szAVCdgBQEi8LJz7Dm6cFXPlV
6LcoUjupzCmOmiJgGSbIm8cNeUmjc7I2sRART0x7wDnejV/yyJdVSGo85gB+ZEGKQvJVc4p+3BAO
ZHyRRj3bvA7zGz6Jw9H7Xjkyjyq0SSBK4Ar9Niz43PMy+CQb1aYtjv4XbfQ2LSG5yKS03U/7/B0v
aPnnQUCI2yGY+TktfXDMgjxKVAhHu+Kz5Q7KvJTfZKshEFN14c+tNoPMIghb/5qro6WlLlVq4wrl
X6HtDqh/c+Wrmx9ml9/5MqQkqbUaIVWRXHSpZBu1vXMr8baxm+4Kh0GvuaF2WamuzYxwB9JxslXh
BqGtS1+uF7fduJSSS3aGGtOCPvCRxdLA/lUGxuo2CKB4OaqryF4+WI03fEBRpIGYMKkaaLXXF5r9
Hm6tcqTWhlOT0jkCkxPdvCZqfWlCF2ucvs77BMAVBRzMVGOPNgTB8VLHeJ6DU3a0YrfIRUgRLpgT
E3ZTTGErZg8zFFfJIy8sUKNsheA5CpCIaes5bwx+bByvfEHnFQeu22SymB71UzkRQSnVCyMXfGNJ
LXZ+/rbuQgq6wCbuJ7Gu2pMRoGqJRzFJtzXsxlNVzbdn/kKrtOa336CRsiRS1JrKu1IREIK8OcYW
yMMkBAcJEqeJ5UvU9sK/R9jRf6GTj9sa27itTY2hUdGdbEGWUCL8faJNLR870m2yRKDNXS1XhYCC
wLYPwecB8CIxN5v0D1IVYqGShqBZiKwqA+iFChwaopfMt9PYuHxbTmKFarrn/ZtrTv4aq1Eh+dOk
Nh6vVIalQ9BkANvNZD7BQI6PJuMMDzk6moauk6z3sn+ch3JKCWpfi6LDqiy5u1YsI7f/hC8apfxO
NuCKXlyb8zYMfOUQDw/SrnkaCmjBJyZcDtMuZU0gss8UPHgAKfec7mEMKDla4wc6vlTXmGfnUd9Q
Z61+zZFPMn6ubW3LWtwEzQ1qUsVeNN9sMtRhInaWnhjbQk0JWW1+4o7mih3w9i5rULBKwHpcuee/
04BB5SJzvm/foQt3uRF6Z8KCMmd1cHdAyttNxavy7Doay0Dtm6AX2IE0DkZRmxL1ZoJDMalSaKiZ
/SaY5RnK3e5kxaPbpsKowng9r98jMJroSRMCwN+vffGmGUD8IiyEOWFEyWj1MyWt0I+qQGjkkmZ+
DHsPyDICMjcxFV+l4l2HGYQoCNplQkChiSQOEVEdc4byCLgih6huOz8eb6/hbfoQyV5sfN3COBGd
m12aWzvGhiN64fDYlsjp6KnKPzcqR46NwuSoLcd0tuQwxqS1Kbqn/AG/QuqBEigL1tQvWwCgrOkE
rc4Cn3JaNvpdEfHQLcJ4//lzay0RECINuN3S1e6fZjRPvMcocbG8TKb9le3cwt4dP4DOwyKsQVoS
1wIX1LCR5vDTbbaWoh36oGJUukm5fCEC68sFjPj4ncvKqllYU6vnHNGokApwIo4Kv4LgA/brdJ6U
erlN3BIBnG9xJLVhuTmMdf6Nvl4GmUESRZKRgsOtk/gJVo25i95CHBcefo6Dv/Gze7KlGP0wc+35
YgzyJwxJpCMHVCI5tFnKgzjWPrXAggnzc2SRSEMOq1HsjHf7X30oLoAn2IVu1pVeSJxA+NjeN9oA
CICxYJxU6AwHwvI7uv2/DHgqtfvcfn6LoEKXf24IZCtBizSWEIYijcraXvAxqnrb8BGGe76VU3dP
8XNnxQlnsGcBFEUPzGntA8bGcf3RG9FLglU3bE6kY5k2hMzN+j2j7dK5HsWmDYykhZN+oh0P+CRU
xZHl6M4SSlLkXaE1wJ4xRm65cO1VvDIpjpE2M2VQCU2Il1e8tBksKqFSZ4aWN7vDGCuZSJADn2lH
n+XFhZ5DhrAJoqWr1WSHGhtWKLnCS4k4tNRSv5AJDP09RYBVhhcsjtJrQ+TUJ+ubF3I7jrPSSsR6
fPTtEavFC/+wH3CaLm6WF5thFPsz/EZtzMmWuYPcFIOMkOnTD4bUVHS40j5n3NKaXKtP6zoFuX57
CkeFNZbeJuFVuQXdyjyry19qhsZvp2gO1gh+8QxubUbYi1lawJCia5zndIsvDAf0QxNioAaF0TNU
1VNtcbcgj4gfV1EezAA4L2mvh3SEiDBOoRr3K2bvuXEnmGVrXVO3DfXJ3hdAAVRYAf0n0AXuASdy
nElaTQZg07WZLY7OaUmqH9NtppQZPbg4D2MdFy6e7I34cTmNxsoMr0c03IbALpbL2QtPoWZrEVUe
+gLtTK3iiTJze5e3ZUNCSPDSdGRlzx4PuJ5q1/CWq4ks2IENOoRA7dLgmODcPr2SNFXzalVpI8Gl
EcxNjxZbVuVZMX54ykhJs1QOKVKx1226kwdArO7CeYlFP75FbBJUvhFCpIfCZx/300TAUZ4RvJfH
nrFABvJvrK0wHqJe3zxGFUH2AXK0wyVdGfecrx3ihyQBeiK+UI1HxHPKq8v3qbplIa8/pBlA1AMd
PGw2qLy3E/HCPaBdRU9zO+nZIT3zN+mnNU33VLBPM9ABrPGiUbQUUZkuh2KWNwD60/iFUTHtTuTF
QIgRaSN6n3oG7lwnGTxTb75kQOvg/FM8EMGohOZVvh4HayVV2jIlDnAqIfh3ZA15mOE8C9/7LP0x
2BAZuEwalGWSudxFFPIA/qcvqy3aMnXFJ5nOF9O2XpY2QAoKwlWOU/+bQI3kIuQlyLI+OaR2/Ruv
fWzkmw4y/ksxs7ckONc66VbuWCsBazfyK5d8rXSYIvSqSwa8T/1Spb2syqH5FcZr2tRCNFunxqp2
STFTNEDg1PGFjZLAKK0eBtZ+8pCbqOuU09Ove429fAx9ETK2ATHrJLzGpgV1n47KI5bOhDGGyQ28
/4ZUpYqaPqwhSB5aNngYEe0dFLHdlILgKX1pHkMGLXKc90DhsdJpt006TR2J6F1C5GHouUMwkqMn
xtwm3mZJxzRwSVrE3TTAr8duQtkg8QY4zpSoieHwep0mTz4tGZpK3XMlSAVBYvBg96u/MZY+y30l
hkdtGuajawgD9UdSCD6FWSCUql8LIYn+p81pW3eXesHpvZGHObQXO28JMtbsDvFFUzddNg32RsL8
TMXR75KUDAjsnRyD4j+poJMpmiaj3aJNoqV34yRzp1bY7EnVyIsOPMe89hiCFxp1I3xlEb8Qltcu
YnZ/GryUHM1xNoEiK7qyefKqsjv3S4oE9x4gFJ1qu+qdfhjup47snukIdw08rbX/PsVvEqBw2V9o
6HijuSK4m3sik2Q/qvgvJ48e3dhgwZNPvUFDeYVuonwkLOMJ+BdWkor15yY7etRkfhBT1xFMYQRg
lHEKfEwIXrChnJBEbT9YmQGogfq9ooVMGbzYreV6Q1srTDso0NeRbP8kg3dlHsRIr8sequZTdZeQ
9b+XuJZtzzsMNiMuf+G6oG4Rs/jNyY3yuCR4x268/xIKkM1gDB0RvA76aLkTnwcj4TR/0gP3EZ16
yugBAs7ze03awRE7fGOr1lAuu5+n+NhX804b3AJA/c26aCACpNn/4C4hFIhweUAylZQtBt7kThAU
uEjMX7YJ4zjZ4c+svCFB0UvABIPwAUAVXTaTqjKE9NEcHNyvty29lpds7JHe26U9ARVMmgujakRA
RsiPnWtToPDXnetodny5XObNZ2pxbnvvaLp/YpwolRviagKCdNAviLJjH4brwVtwWcNovgNpfKHu
L4LXXpj0jvgCtCJUozQrhx2ocHEn1AEhkBYUwa9PAb5VKgVF2S7Q+gz+uqA5WT8DmtiQwmo6N1QP
b7Qi1aZj1a1orY0aO8GWHTUFtHpp0Jgs+oV593nipKH/kGn7uTsapLSDTrcsP+dwRMVRRbp+PzQ2
chYbFY72B5bfKOXjFsbwFU1pNtZVvxBxwH1sqrL725ryVOu9/0WXEL02hi9Hmy9R2FbOpmHPfV90
M+fqNeAgEu4IvWJ/boIxTnPX9ZTXIMy4l8G9uZFDZP0MAmyaRy+lNJbTLkDLRUzpXM15YXjZhweA
sJRf0BwlvsfnhsuWYbvixwKVd9oj+97byQD9pi7v8PYPINiquGQn9GLOYHO3ntOTYi/5VeXPs1x3
ZRhV0ogJ+kSeR6HODxLsII37PXw1dCSdLqQfE75CLdNFVW4d+BwLS4CgM5JBxoohMknXbd2vdFih
DMms6TElpAVGFcpRxqP+CQ9h7oK8d0qtda0AMx2AIM0zDpC+kiuaGpqW/uum0OtUVyxzpLqhrdo0
inX8aTejlq0VgA8aFaV0xn8cCB5oX/0vqKxdwdzm+1PMpBPRvZRbPD8+QAoLf0Vhqqsszsg5+0w9
9jSELw6YtMvR/nHk3slxVTYjeZAatIohUpfE1iMuImLGj14nbI3b1r3mQH4VclDmQzYTORw1kKDH
wJoBaf812x0GeStPfB1DKfUPLMc6oszmBh/rmunUInsMlVDbWr5/GoOmfqKETd/mo4+qzJOh/3oo
qf001RjImUvwOlsNd3LRWXhreLKmIbI4T7KbABEI7m6ueGnG5OfLUz97vaaEYNwvaJ4vlm+utzzH
r0oLsVAn6ze3Mc3um4gjZ7ShtYIMwPbEi/3ttuy9atXW5fw0UUN+PTVjXnyM07LGbaPKzI1I9d+n
xwDh/01XYLZMYqRWN7MlAlFikLc4ai7DYtTpODQhLqq8fl/YZ61imjjmsdZnCOfNqR3ANCTgJkoT
6TocZb5dyzi5RSb2hRLxvEDSg6OLxwwFSjTPccfmX18iUnypZGwN6t5NWEGR6Xl6/fP5wkuZ8xXs
LneiU3hQ4L17K4G1rdPgnbmSsAsLiFC3TosJU12w03Y2VkKFrTsTu4a2nRDPtjAJ0X+7az4sf0Aj
8C+V5ivOCOevOvvTuGaAnL5Wly+zz0DoFvgsRfpJ/0tEpr94FIPyTSi2kVUAGs4vXC7I+M5Gvc7h
1x+xUB2YjAci1083u8Hvhwa3O3FtMhVxaAMMGr020aU/xMQzCPUuLxAzClWv8aREhFrizzQRoSyF
v6gVkyFDFDb+UAs1XYlfEzbdg0Y87+pCx2ZMXWlyXyTlIZTDzI92OdRqudazroricY4IH2fHJ0os
pxyTKpc8hyz7eaO8R61++Ocbsp9rFugRXgeOYwnOY2TysGr2v0RRSql6D1j8xETl8MAObxeZjQ+H
v0JeKSUADAoE3HU5411MvqydWKKBByTBWpsFOB1G8VtrjwFvXApgcDfw7baqZbAmKwoeFuc++0gR
EcKVxL4heQS3Dw/2QTKaU6HAiFfgjoQfA4aZHH1KX5rXzQyQc0OklK0EP//7cR7khs5iY5v7Twni
xXsJFesTYUNl/dhu54uh0uv8fnvsOLDdoidhcbX5CL49NlCRgiGzkPKB3zwNjNttfnPzLZ43NQ8K
PFZ8EOXsmQmH2lINYKbm2Kuwzp/+RB4iQJGL5e6Ugu94w+GPvRM6pNwz1I9NBDX5V4O9KZ1UvfzV
GnYJ4ojhjN5LRbgEK6uA1BzGmFB0tY4zQw5iH4Gd5NXXCCgx6sNzeoskRYd/mstwmi5dhev43sqP
hAdzPzE/BGEeMep3NtVnz/dteMHy+zcs90pdVbNtqRWcDjfUiwlRxoMnlP7M9gl0DHIfaPshYqWf
/aygCnxdvc/OOitRk//GyTGNNWnF3evgVOLng9eMjweBwX9f01KrGTMVQBMcpxS4+SwFLrLLQVTp
9rPKFlZMc5WECxN0y/yLEVwc7k42RM3DWCwM0FYTiRvlFK7j1QKEeci6tV4OUkCBZ6Wlcc2YYRuv
Qw1otrYaT5eG57oa0ww2ZgXS59DwzaRPrrU2DsiE+uuNooBkGEAFaP18PSfPTzeBbNjQQps0aBvA
qpB2b2o7l1ihGzOPbKe72wZHL/oibqru88W1p/oYNW//l7PNcUK5W5Ur4G1TTw0p2PBpfmORvqTG
TBWaTIXVCSOoszWXCs1IHkCmsZv6kyrv3cPWDnmoSfpXsZ0mhas+dKT57yjpvw2zIjZpu2ISXQLU
uRsKj0fKzWoz9pNcbaDwMBC4Avkx9mmTNOklTiq37OOQPvJ4C0PJnsYkpMyZ5KVaOK+yH8KT+GF4
6tTbBO9jS/EM91X6ZbXdijw9Blgd0DisdEuHkwrmauogobJgsbYpHL1l0be8eZhHPMH3qG+UsbrB
IL83UHqeOfBjcS5jxdCbg5J/6hcKmMy92kWy0W2wEhx65h2UEfUn/rqjO/RzXGqm0eWHalkpVZAS
oPNpz+oWfk+9lWXt5F19ahvuVIurtG+23UPVZzdQ3zcDkJDc/X0iQThdHgFWJd8YG7vHjOd5V4n9
k5d9MA/3msmM07+hwZe9Cay3XWUVqkHUfsMxevMH61j8wQHDJnAiRBwYm1QWa6Ha6vuE/AA6U3IJ
YSYgTfCS33dxs1INsNajOUDOtmPfsHCPH3DgArAu6aXP4QIv1jsT5aSJJMwDxJFClE9siSKylmxW
I+DqhNZD+eSoNgtp/aWv+Sfc4MHX34IwYT0kNo/reNPotKK7to829p7YV97znOJtCsn6Hv3a+kYV
sHGG4oDOKsE3DpYLoKM9Ypad6rM4rHz/W5StRQc0LSRazetKKvAV4h17lX9gBtBDyovDkQSxFs/0
kdyWihqNzfqh2dnnpHwZRikcpWi7V3DmUqBiAach5aewnuVFP+EQqN76Ugv80sXnUt+iB9Ma5bQq
lvNpOwDomx1T9eEJPudmkNjp8tzEdDw2CLpLBn4u+iME6M1JWFWLABXsMO4U5Ez7HpdAvmJAHnem
PQhQB/Ar8NhcblJ1nhIEb8ZH9gEwzVn3C+Hka7VtFwjQ5DUA3U9tTavbHq8K9S/VUE7WWVFUUCTS
zp153wOKztmJ4vNLaEMRif7RDgBoFl+UD5T8+NoOelJCyQ1Hp5NZV5PsgmpyfgIGvVoaKxGBUXFc
umLeHUKxhvTscxaEd3/8Sb1ER0JJaxVcq4PFuV53NFqDtF7DJzIdpdNBC83lyyO3rSMNk5mqG8tl
15H1Q284bvrs/Uj9BA3pajIrGvMhxSnziMIRnkGGietzJnfJRWTRe/C11OjoY55emj88MbVMpSxk
sv3vsgBMERENVSFq4NKqY/C06iszhWaEghLUTLbvolQSQ/5QWAMBxM9SFS40AGIEwoNRN0aNiBLm
1GKIxBJuj9VZkxMoxkwcWThXfUDdtBxylcPi0jWY9wbc+3hbDehE1c3fcamfe2vSAzWOZCiMC+ox
uq7CEp/FP83Lknc2S9Lnxu5FrvES9mkgSVpy4KnEHlLBkxGPAn5TnCf6ca/R4klAiFEPVoZuWoUv
akA4rmiMwadDsNiOHM5l0CrIULmbA6cnfQ+3r0+oyVTn6JS4mkD2QSlPaQKGMYCkaIWJGtPwoLYZ
BR2ZOckq+9BYPmwBmBRIGvPCrpLKhv1/Bk11iFJCdD10mZE+aWzAPM7gtO1psVDgO6rhOLRro0Gg
lzVrAOPv/cKcCe85IxEozWQwkAbJupVL7gI41u51yis5i/rQsQIJ4GgJQV3YCAuveBbAgbh+MSry
rHd3usff0DUUsA0VdK6glId/WYkN8tkOEWjKUd3foI3uLFPqwbBwkBG/lw0+iK1q5GgfbzgjtAKf
Z/ucHyYa3wL693DAfjwMlCmsYrSUaBIpifUatbp2a6DkdMGl6jObqSukSBxEIYBUBglMLDsKvRSM
r0uc0UQDBkxZzZtzQW17ep5MSgJQZvsI+m+va31le4rYJZJCIstW2hvWvr7gBZvN7OPkFzWJVa6c
tBgbh/ItcxpHisYPoKr8cU3u/U5zaHYYqp8XMbwShV+mJZIT2Lvxow367lmGLyguJEM2ZleBQ8JK
M2AQWQVZQC8Bth6WQuBg6wWnQ/nJC+f/ehFhp1JQ9MaXxn/AFUjhuDNL+P6+YSNZZBm/l9X5LwM+
jCJr/TGZUHct+AK1Tf/fo0UiZyzvNU5NXpax2NWsAWZNsUO0THaMwOY5EVG7scz/4/R47KMwOSV1
LrR6YS3KWzL2FxXcPv25/m/6SwnohskKyVpgj9AeLIzmjJ2H6cUmEZSCB5XfGVgy+fm474voVndX
nI6XzB6qPc26h1nQ2psBppY04V0wcAd2Zo18YexBpcRcOlPgDURfGm1ZIbpw8kFxVtMLndoDwBtI
VND6Na4gC0y2cXXE1ZCnhYkBej6dy5BlIpX1PKZ4fM0Mpzz4GI/RlO25whev9w+O7pj/RvXaoJtX
PDOBLttyRZLOL+SvTGg6omXSzPLkbNffgFymcLe+G+5zldoa61pBi/S+egUC++jHcQqd3RTmE6jx
/guzS4+iikK82RIK8qjsRKIbl+7ClyBukI2ODhGE42QFJfFb6TZVqKJH9ucB2Tk2T73UYeE3oedO
2VGH8MXM3rbCJWkhmDZSmKc80/gkouFzNxl8eP2ELHlqviSN+8ISBSvZNCTKadv3gy2RwDXtwiD6
3Z0Y7XMJps6nAKkCo87Dgi60H04sG/FRHygPeYISndZQ6jXsUJ51wmafIZjLvp2Ubqhs+A6Q/cAN
5s/NRfKGqE2b5Z52SBini9fc6Mgs9Yr9kXvY57iE+A3SHH/BSDOpNl9Eo4zaij/EaQVZCMt9O20Y
u3zALgUvAeLtGMgOb16Io8uHh+SDU18kRHpCTwyIrYV/wvJjwPdoLK/z+9It8b7xh1/FpH/gTqmA
Tn7MDm/jESAaDGpGLAxW0fIPScUIvzFAJX3R2p9Rd1V6a+YwDpCFjRTq5QSfjeXmlPv6XyDQAh1U
OU+WdNTxXOAfOR4tqBZuRK7eXbEsQEAbJKSlCR/eUTgIbosgekHh/OoPTyk5MtYRMK1naFde6jyk
IhBqYQ0hIKKwyLy4QtdGbrbIV66cCSVeMZDbx5Amhx7u0saJ3tGSZk+MrFc1JD7nu+caWpWmDXk8
Wb5tb0uMQxI56uqnkKJotdl1QRvpmgyrEclhfvytFAdPfpI42vuWGRyU7qv0efkJpQoSwIuHga7m
FoKyu41ZLJ5Nw0oYa3lqaE9ms6Y/Exlf03szMDPCFbt9LyUSeWJ279hziDhwx8G10ezc/CbLDYcA
ivHTzJUzLnkxukO+jky0U24Atmj1CCipl3a1L13r8qdw30W9fSV+gC8xTJQZgRNjAkXIA0P60n6N
ZQtRLFHQNXQgsXwpJH6ReJjqLD800wEbNNgw8NtLUpC4f1bu4EoT6IUYXfbBSkiLAUoHXT3+3Rky
ktChHR03QawIAE5o1HsvITUJ3moOO8MMLFLUjCPeoFtmo6W9deA72CFvmWpyYMLJIiiPsCaB3PPJ
+3wXDx8L7iuymwScck/MncyOlFPyUY616/Y5RBafVJ7sIwic31WUtWP3iXCDK0r3/GY7DbH3JIxR
igIZNVNs26U0bhr1EfJj54v2SRjQZ2lQc5ODJJ/MQR1j0AihpFJX7L4sugWTVotAGrwOf9HIu2lh
wg+pcUMcW0k4XD7HnMaIS/ZQ77qgUWM0l6/xh9DaWFCGZOlegGNLfb1WAeXHQOjo6IqoNZgkwHL/
a3DS4rTpUgXeGw5CTbTa/VNcMutgzgNO+XHbDNljoj6KcupxFn6XZrx8yKwmop25xznimAxjM4dd
Tg9BjuToaDH24LBwd/XL6QDdfNy6FKFmJLJ+MIvuKFTfUGvtuAPvnS18nm7zw0ID3ECnpnySUmH0
3LQLAUtkfanSmPXRCf4qsF8mb5vLbeKvMbn51U+tnG27/a7lpzKkUC+TbOZSFUaDYm4khSkhxrXP
dTxqHklwYldWEOobGjRTakvfeO54JtE5bkiMP+k7XNxJPpuLjvy/bdVRqk7J4MRAZY7wNKLX1TSz
JiuLEj/9bpCLwbrj5YZ7vM/ysyCCzAX7iknCoqP4vdnnWjT/SAhVGbqe3saM/yH0hq2tB8Ge9hXg
YyK+HQQ76inNUM6U/7QY2y9JcnkJpyCfheBcHte4e+zJX1ZCWAic0lLBTYw2f+D2etImRC2mTfTr
1oNgmTOHrV7S2u7gpxR/tr/NnBiVUypnnKMTpHRrt7bqmRopbnBPdyR9XsGV0NZFPJGSbOkBRPI+
9J4FMWJz2k3tqJWTmWsJSRLj+2RH+xyUAUzdoBGo6ZdKq3xJNjcg4O40IdFpGa7tNHIfaqRDXZSw
mDZtUu5geACeTJxGZONwE91yAzYTqHPCMN/XL2mz6PGtvWSxee0mON5Kx3kwPhJ7auiu5yqgZAf8
87H9GDIk4k5cAg4KLSg/4vu9wkq/FIcXn78MICjD2q4p2MqgRj0DP2kJPqMoTnXz3yTjL9/9zWLz
7YIfkZjf5iX85pltbIIv5NvLNUoyELk+UFPMxwp7Rq05dk7oinoly835f56ugEi82XdajikjPOvp
oM5ddBjSmkyjRGhjGKaw/jdbXbWijhGc+cinQl4zQFmBqFi3Ogpwfh+AVfABttiSXET2I3SZBzOk
/L6EznZxT2bobLj+3+eSYuhUmoVv8t+3lssUSo0pj1/NhqtvXu+2M53NVz+G+qOODItr5EFRu3XN
W4+ACB03odrsbgqL83lrac6W9Kj6tkbKsDaKZ6DkYR5zhOMzUs2nIAmYdgC4Qon8cZvHGVc2VmCd
7iNx6lyctSopmN4pbFhRqsH1X4/Nfh1IjDYibIxft6Xvh/4kBBAQrIyZfWBBIhOnQSMR/aXFVGXR
4yo2jyCJMorABTpUOIfIhNAicUIcGrKd9bgXBZmgU9bdNo27cqWbt2UCAHOtRAv201SauZRKmxVU
NKuOcZL2y4AgIDg6ekEDqBkKXI66gKzY6DrsxcTIoiYndODQH4zfT8PISZ9nQa6y84nLFMDczVqI
qUDxcORTqg6gEeG2pzmZu37Mdb1GKX2zVxCmBtgqldjd9kbeLUiiIUrcpYtBN/I7i/7SONbEGfdJ
aIP6Df39DgCEOeTDhXkJlJL8DIsyOG9spG3bH52+Zlye/SHLn9EKwmVtJ7X648UPMk5taWOjFEz+
8/9xJKaVIVOKOgDJME/6R7r84Br30K7jOVD2yvh3RoRyM5BNfx2NU7nUpXdS3vbgr6dbsRznKmjF
AAzbbk5nmE2LUM1rfehXqF/y8YZjThf82FlnpPacSwNFuDiRCBRx+IIMeuDguH93fuu2UTj7WrtD
yoVkjOpSgyDoVBdrGXGD0mSnG0fZ4umbF+7vc/hvHDGHH+0B01Q9odSs/PUqKYsp0OyC+nmm9igA
Bg5txXmDydfts6rcmfkfFDlnRin7Vw6p8nOZIneLMMsyzpkd8K1suRdhFMrWbSW7s1DfPokuG/QW
ObGXpPoc1mJDR+DaAdERpOVeUgGUrB4CxvyeXLh5MNFYmXJcnNQahPl6LP54axj7CmbAOkUZjiZF
aeXv0FKrQMHbcWpX5wMiE89tLYynxrc2proHNiICPy7v5RBVGBlPoRnV6QgkpmmJHHuUGY3fUWPg
o9jqZ7TvnfQCnyoX33RZE3oqkqIhtl7LlV7lc9DtQEaMZegArhUr4lG63MBKMF5Jf9a1FvjVV4aW
5J36aIRR/D9/nyzKaLtrOBqpeAtqhYsYwKxu2XgFwunIY1vTRz83GkH2HmwYWxrwKX7nJh3EGRqM
KsmHsHr/00qmaWZEZAF3RyPvCW2lJMpHbAD2oSbQbALc7WhwiJpTip2vsA+n+m6l/36NuqxEhGOc
rXxBYHaj947N9ItlgecIwqCnBy/sVl8/+z7Di4SZSbrkzktzHq4ml/0+EGE65LjGMN717qit00Ja
BhRLvxdoe1H6nPrF5PFiP4OxQT1eKtF4LP/KeQtPrNRBPFAUSz0aewldb3vWnuMnobE0nOpSzSXB
mdMeO60Zz0+9+5ITS8Ip4yWx1xIGUcNDSmZbJtjFlNMGcijsXqckqGU/Jx2F6VSo0yqLavEakVlo
VCtT+EpNglHXt8Pz324/0rm48/2KuqiQuxUG6GqAX8dm9cueMUL6mXAqs0AzLrItviLOEtux7EX7
b78vBzbNzsf8xr3U7QynAatuwuugYMhAiH0+hoj7SUgKS0UwVnzr7MnwuqGKbmjGX5ApyPUeg3iV
Y30uwsB21S8/XM6+Xsmdv+XoA/RXShQBioSkpLQsNZ0LF1X9uca9idxyUOuLVRqxA82TJkBwHscc
1JYzmwhAJ0QYINcoX2ZGt1lmYABPXbk2/nxmRNsoW33mYQ0q6kK/SDb1/4F2rQCbDOtyM2+tfLPw
b7KW0trsq6y+6PEKtxke54fHed9wGW3q5q5y4nqhv6RjrNdGV/6PSODfOH6FK2VV/BRgX7/dMgf2
/Vx/Fvvus/hirVjcAG6VB1kAE70NiLMfjSjJO0+08KsuJd4F+uv5eZ8ArXaeWq3tdIiA3lqQfOAH
any+bTSZVWzenAOC1IXkAmj44Y7ZJWhaWoLRfjXPyPq5Ckt+H4yOeW5yK6Orh7PikykAaAffrcbg
x5hjW5O1tXO6Hcpwat5ekqbhP/52Y6JvS/yz8d043PTiXXJnMYgkSYIqnEpSoRrDIcuSkEL4oJwH
EuY2EIScG78sLM1Q6n2GlqAMrf8AsTmLnAXu+fLrGkpioQrd0sFBpnr0elXPdQIzmqAEInAwaUX4
Id6LdZgvxTiHD+m8zYd6wUGrRkLD0RsKDDs2N3phGjtFX4BZvu8efg4qAUSxViYruvdNYcFkegnr
zALVFczGwPXB5AqTSNCpds0STXY0m4N63ahcO4CZmwjHZ/u6478LAOB9D8JMj7vRwFGS2Lm9LZ3u
8KarPwF2UHIHvLOcownB+TwNKReGgYJ0BpQYIIYxLls7moALsr1ULzHJl3uI0BJMgYIvHLMI5xFE
n462086TDcGxuOc4JeZDsiim25vt3crwwBxe35Wrl0caMTkY4ct41eE2eHYAjQRzHM1izADvKWSu
suYa82LNHgvtD8zi37VM3M3jTuS5i21p5kkb2B2lVBhbe2Rn/RyIsEf6Ac/xjsYleoz+wiX4490k
HG0cAPSX7r+Z4osHgp7DhXpv7XEMOFJyCBysR42bQ2Hu8aRDtNcNkmCVPzKKyTwC7IEwmF20v6BW
GPSVRkncyby6PPkmo1ktcv2B+ZYWY/SMWwTabmoQi2ww8Y60d8q9W7d6Wt9u+9fkj4yiyIUGZ0+2
r+k0AVIcKqD7Z+o0mhDq1oyfVvMSIJZkwZ1ub9NTZMj0weM1KGqr7I215pbi28U60yncv+y4XR8X
2h12slQzTTWlJvBA9jcAQ4HuRhWAAew4z49DX2sGkgQ//FWoNY2ZaM7feNwMMu+IQayISUtM4wOZ
gzb2D9vhah/bRjcY5/c8KF7RcorKObZG/PmugHfflXIvN9d3WC7zYzZycuJCvxQ8nOnCuKwOO43O
qUVoC1qXzH9x9wu58h4p4YZvfUJ5RrNK5Ckawl/Vu/i0BFDwQYelZw454e7kn37pGepxIvyxykes
Z00oub6REVsR91fq7AWMfPFvCE/luvIzyk7eCG9cPW2NP1klEtXdMqC7eChgTBflIyLjNr4ykMg4
7HnFBJm3K1jNhjJbrs2Sa6PPsoVJsVrnmhrua45wT8CGMZIXENp9UHzXHx/eFHRPb1RXyZe6VxK+
BntGmkpP/7muUOGdvdj0CtpAFvksMKTdgpJ2nOG+GI5mkhL3LlSwfsch9q2Mr82trTNXnaXbWo1B
N/oAq8jhcxitDjZvC8y2vAHE5Yn1ZnX4vSo/HRYY/PBFMWPqu848s5MrdKnDVA+Sd10DTeYoQu1d
COUHlm5HpG2z+tEd565zGRzUPKJr2im16NJpKIS+iqvCyeWBurOlpCqikdEAhdoVVs1kbVXHKnsD
5u8uBGfXGrihb3IGBl813+hsP89x6mEGj+T9CL1fa3EnCFRc8p0hGwEwQHLFHgWOGjsYm4gavM6q
ilebuxkYdM0HKnwtFlu5+pWdwor14MGXUhLtmuVblfgI6DgatU/ZoHKLKx7+xsmWHrVkQ+j/NBfu
73sbpQif1IE0n22DxXswIJbv6x+r1obEpETR/j3igO84Dch+s2nyS2fkTJhihn2beCZo/D3rpUBt
4S7ex9cdwB451GWim9U1YrK80PVexIPpxv+bzJ4PcU9B00Pe+nAGH9Bv/SPEktrRlN9jppGq6Sf2
64I7uae1Dzq5bTU9N1HlTho6KaIQZ9NLTjG+v/iz67RLeL52khAuBF5PUTNa1RBQmeLh8TtMrC4z
lBhnf+DKOaswQnyteSahFHmsUoQJ6O7/Hja/Kin5VrUJy3edSWEX0xY2R+KZEybftV8mL+IjAbQH
F/tXRPaxafwmKOquwZjncxKPzZdyH1lcLQKuVZltdS0IWjJBZIJv4SU+4byeDCaPydnwcdcu5CAs
PBtaNf/05E0yskGQ2Ra76HqL6kSFkYDrWHRpv39Lf6B22DzyV33eXYumSYIGjJWkobzl5+g4YN3z
e6opRw6MbRxH+OZd/7cF13Ui+Z1RPe2KaHS4TZ/kE9lbBpRIJePYot/nT/U+mDn/QEUri4QcVcg6
ElcYZNULEKkOJGPsySYQq5L9HFuEhAjqLIPqopcazrL2xn0ZH1K/j52PJDl/W/ZcPzcuoY1Ug5vV
EMSa9bHpfmq8MfSQ4bB/e4qh+ZMJbj7ip4YyzywnGqkm3rnKTodE4spLTm90LWD8QIAg6PtvXA9q
98Z6dUUpSR+/QNjkwRQ3Lum/U46JSz4LkKXvUMt1I+cNy18KioFkeC0uUG4tl5hQYPLXxSLZxHrN
oNn0IPpLTXCBMnYdIX98eZ4+pgMvl02tTWVpZcncSsGAlIGSfc/b1FUtZ4+3PZKeE7MTzB7Npc5G
UMqdNRUWgImqTt7fxu9WBiRCNs5xNdFqMMhbZ3cwFU5SwfxxReJdfZz0jfWtwO32v7e6pBifZWS7
8cimB5ZUacXDNiA2zAeMmmnmUn2S6kLGu345HFo28WmVzDtKjndeU2xrv8+/YQELo1TyhZay0p3A
Dbm0r5OfvMf4fJa3hCzA+IIzxNwi8ZF9tbDnvyX9Xmg3vvrUpyeabgEQ8OmlM/05Fpt2kXSzzUTE
f/24SGyOQZD8GPNXK28T5nAReU7/iqX4iQ+IGarpUX9d/ZvNhAz9E0gvEVF3zeOybw1ltOUe+wRI
Ob1Po7OMmJhzyJcEGS9Bjc2hu+q5pusMCDruRjdaxXWa5VpoZNTWZmZc++LDgh/trkPiGMXJmviM
haOMhlFpJZ38O79m6mKjGNbVhMld0kExsdJWQ0gsED4a3Iu5HHd9KXttoTtJUZbY0MdttXDOwAOe
zcsZuTwlDutjWay2ixJpduihWWDzu/Sx+OORYU2IZ0MeOkUHaYXyvQBwW0M6bEAbgcLr1wNObqhY
VAqjk7vGbMKeODwQiGo0+YTCWGyFj22YCj0g75eq5gtyNJpN5oMkmXrI+ktEpTHFEvadP+UnL0V4
zgie3EgeyxoT8jGasxQGdP1whdL9e32cc2gTJCigUoVQovUfQY++XbvcBnLXk+v5l6dDODJ2VwuY
GZw4QYcc4NADfs6817lgST7FI13qJrbG6htAkZHxY602P4mO+dyBr9+dVF9TxbA6R7CxaiAYxz6Q
KsAGQeOJdoyC7E6tOM/Ijie82LYcGhMnm7ztRL9mXv331f2tsDHVQhvxCEF/N454nRlcXPc4T5iG
/BCLRe0UXQS3m2/ReGX8Uw4P+iETrnnsTn/jxgg56+E8KqRaKUWGV9hyuTJsEqgurR+mCNlZnZHM
2B16ZMgNuJiMMrm36f8CWhQTSKUMQEXaP7qc6VABBxQZsGyP6L5rYKAp7zzHE5qyjU63FiQXaKVQ
AfbSqGmhnrmlOoB5OSHN2XcRcS+1FFnsX/EbQDwAR/mhsP3Cnaw8S6zwVtjLqFh/41F154i8a1qf
sViOA87qkApFu+BpVRWLZZ0ZHrJu591yGvg6XO/dQdZzCY+u0qwCun7i9uhX7AF9+zjm5wjcv9Mf
9DD7FrZoOBQQkU5Qa0nUsESFATT2qn6+l49R5kWKxReJVnaRmz18XdgJiDEmbeZ6s8qMF0XHDJd4
EpFUWpj/itlvRD2xosKHGis4kDphZDZYUjbXnx2+/zTbj3SQ92zXKXhmYTa0A17OgdS2IngQUcnI
QJyaEK7z8zaTRs3TchlMsFloGP/bI5aOT4zr2uUu3kDWDbvEc9R6KGC5wBVNeIsPcz64ZuvteU/X
70dbFsIeBZ+7Fj1W/l4zOJfKCYrGMUatpDi44+bowtfitxuoTio8UmxPxwq5G5DTUo7VE1n3jzEQ
Slm1ETthK/CJ3uAVxAmh6J1JrVyuE38BZiUjmUM87e5SRk9sJ9go2AZyDZ9hGXa/IrtzUulxB1Bq
RoYtYKoAl8AK6ywmN3iEQU8XdjT7JGGBjOySCWjTPDd0kwr72dHBhlfas9vOxSDOh2t1/yoVbFdU
itXhZWlTrULkS50xyyo01u1SDz5YCZmaBm91CJVjR28G+5fnaaYtxgaftcnKQ44gPg8+9qclRSX3
3WOGbc1x5VFpXqtYHki3/7UhfYSpwarUPlSH5Z8LwPdKV3hL4+qVxXq73Z4oAIyvkvjD6SK/sHcr
zf34laN1S+tGpudamtt/lWko4Ia6ERBHPwI6A+Ans2JsZ2zEUq1qcdum9xb6kOOyB/TxXr14koFG
MHN13uqXSODf4O63xaSdrlLh+9hhdvcKt8FhsgKcXJq5FV7Yz+4UGi093NvM/aYyv0D4LoVrTEnD
6qB9RmD19qTUS1CmT2qurV34AZNX46RD6RO5znEst1CAa7WxsxWgGLwmcVDBFq2adPlVGSxw+O0r
l6eGuzniMwxjo2/QNB+CNmp0Vk7FrzI/BHo0V7xLWorcXAAW7JsNpOTxvxshlxElSmql3jAK3Z1g
5ifAkY1O8qoFat841obqLmeuyywyfazMYqVxKyCCAY4htSq2dCVoqZvtgosEqtBXOksu1UFp8+fM
Tp+BIQ5C2c6YAQ7H00XNhSV29eTC/xlf6rmwg9SqAWfbdNUWmRCTStaEUK1GCkPIyR63HFRy+KMy
JA4Jv0brwlEQYrDTbPNmiD504LSx7JS6nIhI0VgiT95WlO1wO4lr1MK4IkB0HQsA6BULavCIXyMd
glXpXoxkh5o4MkKEMtVg19udYhxfeaEcFD0SlL/k/3as1JcioW1Yy4QE3np9SDptJ12AkzOYFMfL
l/RJ8XS8kFZMkSRuArZPjczDANVf8UInJISGad3ncvXLzoN52QwNPIBVNszWL4fsEdFZt3t9cdW8
wNzmOx5ST2J6+p69Q3IbU1J+ZvKdVbXV4n2gFoXJB05LXbZmRQtt2t/FKnaMR/bLzj/om9TpP/mn
PKQRQxk3c2mQkYtoKu5D2mpBaAvD4LNq+ObB9QnxcYXU2eA0v3gq4oiqCQ486CN00TYihPcGISaT
wrNgcnpGpZcg+6D7JHg/WO5XfawRJiwlq/98QRJiFFVKBi+rOaCfhaMGlumfXspB9HnPMmd9VLsZ
HEQEfVaAZxba7fBkQvJU99nK1iqzNtq/F1Wj0DPISAuDA3wINMFvAK7NIxYM1RpBaCEgecK7tSkx
3ILCE7MOa4M4Dwb41mL7lJHRtT2LHQCM7OrfuMxQc92ZUtO7tiCdWhmCwe7cEgYNT0lWiJyxTI2U
dW21uxgp1lYFHz6mcnPrnbf4WjAo8tpArJRFGWTV0qmFWa15be8hYMbYl5bgdteUb9kYyapb8jVm
JTzH3IMy9i4KU07l0SfZGBBbWJgocEAXUjHjdgqI1qtKxruy/7J4QoS8V8P5cyFQhSgfVDvglGJl
J3BCojoH8v0p3vPCpjqDx98HSbKctvncxVpaVlRLeCsnmhIQQsPw+EstgkcN9DpskEWsXJLL1Zfs
G2M1P+FsITNud9e5gqAnBDL9O0hdeSk/9kYuv5ZogvG/aawYvEj6C27Ba5Tr8lmRSS79d23CdRG0
knqV6r+izeVzcJfg4GNj7zS4KnFl0p1qwbj8AVjY/hlW0q9jI1K4FMYkw3fi5a2J6ES+s+DuVCnG
8Ooc89I7tMXabIGQwuBD9TTM2FDNV3Ny5W9Bdp/SgTnwM7hoBxIao+wTtNKZHUtiKp2CU8t1msQ9
YlTUgjPuYc8eHPg8aUlhk0oXJjlQbQXTi6zuCZq1+KwT2973cN0h5eF2mHd30lAEsDauTl3Cqv0j
zT49NMVNrDrFP3n/Q2m2DJAtzM3UY7CtZobN0je70Hm6zYOIWW8OXQlq9MAhva0hTLmVbZUh7fOt
fiPMtPGRtV34MMrJZ1tH9ZaD6rAfrvj3kypb7W5X4VpxTnjsfRBSVUP2pcufV+jEhTnUe5Zzmc6q
IiXtRJeBkVW51kVMd9aoC0wRw+4pI+AQtVluBCouelI+/M6k2SOi0hjkthVIHWV4y6aIINxkguzl
YtBMvmCqJjFm5gGUAvUi+FQOlWxfx5ntcVZGIiArENUX4zKU7wDrnWwIJKAPY7azpbLI0dYrhLJR
t356deZQNBbSgOtg7c1XdFIJ+E4eUWDGdWXs1wAtSwmdhSx2pBG9WOw6qdT+lS56pCwfEUp4DvIB
HpbbQUeYy5rSCrzIbeScovs8w5xpbEqLFbPCUIR2IhFKvFs1p0he5gf/ql41MG6ilAsAK3AIJQ5U
KHV7xRpByjNPRnSObGmuuqsJBJeR6tzD/gyShOcKmWOZ+MAkpiLSzy7cdV7p8o3WDpqpTb4q1h8G
MkEHRvbdITGaRxrKj1RQrd1OuTBqXNPeRymJ55wQfe9F3kZZZYAUGB9kEww/dK9oKaovdZuXyABQ
iWhtfIH25Q/ueoX5wUUVPcTn3PUm7scostRiiv+pDMb7ULy9EQ5aTV2aCQMAjRwj20bKTW1dHfR8
gBvwCqXUQsI+gwnz62gd5enwf8TCmLLfEFUbiJ6AM2t72kFGCgCOBxoyuWIMebuIfnQH3hg/KHJR
i5rGJ36TlPt5qTFAyn9BFT2LtaDWRxU5h9jQ0kBjgEfb/k82J2hZafKlo2+fBjlhw83izaXLQAnS
PiIJ0uLrVbfmuB9yxu7q1OL/JJ/BIbkDoaRcGC9kIW9yi1PvP46XJV+GQbxFRYoUXdDfgigOGOA7
UXVyA13nimh2v8jT0u5pvPCNWKv/eHALhHYo4VKyHErqt0j2fqVAUmdnRteLdG+j1R1NRDTBRzV+
/cwDsxKytasULt0Kfl5CA2qOMP5QeQbOpe+nR+ijXm8jmCS1O6gKCM6GNQ/xEpS+AEfSepHGSQmT
1Y6+3ptfz3l9T+CPohh49iCRD9UZOeVLL88s/RRKiNNS5Iz9H+eAqcZOTumwYjBKJ5gl31ClmZ/2
+LjKHheXySgTbLc0dEbB3g8hay+8iq0XErM3nenjB272MfklRrB/miZT+8qe1028sGYOygnowB2t
2jMSH2oLQyPUvbeSPxXS3KJTPa0KDNvSZZjiSwZkAg0yQ6B+OCWTEA7T9LLcEdL5T7WVIoSfTz9s
3yzEUpAcY3n7hehX3A5d93s9TW0GgvvhBh17EWG/g68eq60AQCqVF8htbiph8niRmTmB9Z37IgPh
lZE7o9OZ5lpEsTQvXXvPJz3OOLTO5w0PoWUfFoY4BeXwbiiNkQ3nml+BFVJiV7iuWXrR4jDJuTGg
Up7h4U+TmNdr+XIoDfSkLBklNVn2dNk/ZZEc0E10eigTy8nc2iybCixDjn2POtRSTY/IrG9+fXG9
f6eTuu2uU55o9JGR/2VUHMhJuLSN3SrXvOsocBMjAp6V5rkPfChr2uBcYCv5Gqxel39QcQibmNXe
6eCLIJX4fPqT1BIflWQ+3dkboj/7YIyBmnekVTthlJSGWR95+LfufztS6VOQ/TUYzo1xwsG2EZm0
hfxwhRKCm2T2k3hA9SarO8vHvhr/yersE3Rd2GTClk5942ttCXyXpHxUFZcVIX2uMglTkPKhTwcA
a9MDm/hQZirPNH7ODNYN2k8nU7bbL0BNtiSuNYcQhpnxy2dF12x2Tn3OVaij2Ip9HkIphYXSIONK
n9oC7dcCfciswv+nSzxqaZL6ZUGznI0Kr+M/McR0EY6n/Iwnkx3tfPM2GVBE97ArpQpgyXx3ZV0x
a0cdFD0AnDTvInTCYBassQ49aaLm6619TTytGZXDvwzWz1KytyhvJaKQggbc2CBxWj7yrzVYxYB9
Tp6nixbfCyJrlxbgwckXFMtqmdV246Q+QcgKby6Ii6KjiAVjO43U6X397Mjl56lmYSoNev2LKx6j
dB5GO+StG1PlXcKCDlF7M9hfcoK/DugCSMxF5rL4hhj+tkNW9ajq9AFGImkrkYFD1uUJB0j8qZmU
G8xSGb0kYqhAs+WbcAHXa31NqWcaxLxdmMWN7f45mNyRjleaSHMn6vAe61OSzYoJZf39MbdN0H2x
++SwgutLfAjeciy6M8FQVmsCB69R/16dW3ywccImfd97EIYl0RcttWan8zIMimJQEKp0+YqOUz81
NHR4yBqcF8l/oj6gGyw17E2HLJ4vcNU/RxrCE1Jk0BVRbF9p5bi7J6c+5q9Kty0af2c8XONN0FRS
Ja0LZxQdB/Gsq/ZDD7ZtoIGpeKNrAA7fuKZTQ+QEYpfQP0jJnVm2n72mjBseN51d5FjQqQIrAJEO
zZZhjRtKVIY9MGqD9g0fBv7FpaaY8ks6Nh7kPhKb6gAOu6rkhOAYM968PEGwEDZkx08SS1M3Cz9Y
NXqjzBMVodQ+pUL6QBz+1la1KCREN0bU4BYOSeYrXXaS9sBXB5+TglWnhxwjN7/v+G1vOdGbFley
/VqzGzw5a+0wehk6AI4W/KkfG612k9e4y2ajz7uQzZIgjxMdsr7quczYDErB4c7A6zLmYZr0ml2r
7eNp36JNSDoIt4LcfUngEdR6nljgoLoV5HUiBa32La+CmDqwdO+sVfkwXygN6h2EMYkyUZ8UdrcQ
uN2hSc8Bk/7tef57TaUBc1fN9xBxsI/Hu4LhacR504GcQNiH0e2bipD7+N+AcLraS/rGmR+yEow0
q7k+GA/WT5ATeEEeBwt1vgK9Vpw6EVqyoOi1JK3wTwOfEuc1ELqS45+jTTY+hOC/rYI2gkhlGgT7
C5cJthDSmMftrs5UUBaXYPoKmwm4Z4p6HstEC8ZWkSDYRGCwgIF5SNzqOTMca5ujbX9Yrv6wOhhG
ITUmamA44wRHJ7V/Detns9gb9zp8/EaeUBKa8+GCADSxx1Sfi80h/24L3le0icfq7v/mqXoiZGbL
hwZPISUC63pDDabn1E3kULwXARP2yBZvyoIMHUjLHK7V/KCxSo2/zBYNFDxxwPSMXUkNPs4A1eom
wbU2gEUkDMhOQGA3fYOjUPu9EVFhPofg2+6+tFFPJp1+5qP7QI15lCY95F+MdXJfIr88gpOLWWlm
JuNcnxANqyMd3nehCCMbMPNR8DLzNF/cxA83HIEXXQofobVgMmQQ8s/6vR6wrsBO3if4gGVGc5Md
w8AwOW3xzPmoTPKHbAwPd2XJ6ntATJpr+qX8ASEclX6D3pUVU8VC/WeIV0TSVECBB9oUGjh5sn+p
c/UnF67/6LqQsiisOLdOOPPI3MiIPoDSopgLR9TjsnNxwGSC/ASk4+cxjrK3e1x/QoWlirl3Q5u+
vV97HzYlFJvb79MquabUIfH17Kq3yrQVRZ+EnjIXiu0fpmRBuQbDco9Ko78041xtm8xXPMnUwpFe
xpROQugvoLbsMnXOSeunzTyb9tkgLkLA2TVdXRXvUBGUtdeeaohk66JNATXi4vMMsqybLdGumMcD
SO74YF8E76s8Dkd9uDWMmBn/FNBX7Lar6FWVPSGdcO6kec8pteSkt1+dpWl0ndPETwL96RscswEE
J1p+bYTLkdRCvKVVRx7iD3dcYWvh0Arahs64GyFxp06SN4p7WApIgPSsmrUM3tlWBqhcKPDJIepI
+A0UfP/DNs8P/IwLPkkzAYGjy9V51r9+d0ITsvSVHxBHvt451OUUv1640j5JXbHolb8MW371E4uu
npMU6lIWzZ+6YYd35SOyMDpxHcrbAoEi0bEQzNHJn6vUv8itDwJPRElep7eoya5UX9zu+B8+IO2R
gKpfmcrMp8RcrO1V50dzf26uCPkkzfg4bu+ty8f7H/3XstsNfFUb43uJ/JZyB42kSHzslz3mLjRS
co0i4nxA/F0PHmfn4pcMUFq0pGoBasfTLBa7CMthMbW/0Ape5p6euESGbAuVkpmbFR/Qph0SQy0+
lWf/CNysNKhWAR6LlM2C5UEAsH1CBusP2qPMGXB/jf7PVloD/NJc6Ltd5RMRJH7m5KsdpmvgX7Oo
DMhHRgBXLpznzmU0w2S+1Sv1TNhaitCJT/vouvw+UibtlZIbaSBv18r53JjE7rBJW66HLne4l5JG
d9NCh15YyJaEuq94ayxb4zF3Tx53+FxmoOVo1OP47c47M8aUW5DAalXxfnlLjWJ9cBrUf5/k0tPq
DHGzhLPCgGMGVAsTZjlLcY6v2E01FSKvhTr5ruQFkqfteecyxweqreP30okRoVIr+LNMdE2zR/Mn
R4oyc6+9cnRVPIY+bXBfdWwu/5lmXXmPdjGLSMIX+tXaCBOVqfuF2nfWrskH3ZlUUKN2VNGAZSaC
3497DwTjpyadjXRhPF8iGEU+JRpfszm1jBihEVLVv2EP/0Ciu2/8kc8yLqABmCAiz0a8PNZoB1T/
Axk/V17HpX5VneOXhqhKdCmRWLg9yeraAMXlaKSqRlGwpeQczeQFjRF2ZMRHE4WM3szDeo0aXLeo
T1ZuJDXt1kp6Cd2cF5XmX00yQO2Nv3EcjjbEZ0nVEZm9WvnGOCUbVjLVbPzNPYNGdgn1Ie6YDoJw
TJ8NmIXZQx+3ytbH13F7j9Zw+MTAbyEENf6UN6FD5RsvGN7sNFTDIkOaI7msbIxExfsq/c8cUIvU
8lZKixhJWH3frtzGV/oq3esr7xmt6zHfx67gLZStfP1KarRucA7LJVMh0G3Lad/mknYuEevgvrZ8
/BiVxWKg36C95VIqdXWXr+yUXvjja+fVp5nlj2Qzi47rS0y9TKVOeE1k9+bSmAmmJgsL9+FPAc7r
FKa25pCudKxiRwppz5d78e9pmirELg2wcYAervDx+YPKCtao4V1o4pwd264DTCe9ZOj0FddZ2ST3
pLIj+z0jMirCcWNmUnNlmc2Ky75vBhEynKgyebaX4mDjMtHN52qzwIBml9A9OH6HSaywd/UrGolj
r/YuJUV+vp4nVrCOUYgskB9jfoVuQudfUjRWxheXBEf2ZsweypZ2Exj/6Yg2WQyh6lKK1PVHqArz
3DaNaMYh0Hekjh9KYzxsEd0IreU+Nu6G01yNH07UFy2e4fRrLseDaOH3YwaxWzBjgOcRLY6YeEWW
9ofBEOtTN2JRacZPJkl+wFDnSyohuhQAb9fjUusZQIUXIbyweFdggIr7gPpzwZutG30O6LDD8izN
Bo0oT9OVn1PtP+onQvmlIRsViy8VCnd3PlmaBf5HRCWQLRXDo1Z+KqzSyDDwgmHjjr1EzaSn1Ux9
OTerdAI+W6Mn54jj3MaeTVP6wlrIBN3fSWAMZt0k0uToYmUFIiDQcDmyywSmax6abq0BC1w4YHtN
JKXF0b/T5P1OfWVxokk3Oay+/IgKAOKJggNQ9ZLbmhvX0Nd1ZdCGA3vnsIxbghwDO/eLX7qyIN0i
yXuG2RCovK+xsKdl89Pgb/3FmO5FhRy0moCV0wRGqmRGjz4fpj+7DDrvJEGd+rzzwTgeSByLiK6Z
JLmD4O0vZvx5VTkouTIAqMy9FO52xQGMIahnG/DJt7nD1f49pCWt1JBw52wEydH6YhAlEkg7PQt9
jWk1ctSx5XYe1pNeh217uNipgTvtNbWHRsU+xq/VZxz3LecIC1Tlfor5tM25vp4VqfJsSJ1VRWSH
YAwXIjyilDfV0e61X40jYOwAwbYx4DvpOgaNTjK0grBVLT+OpzSSMZ/QyaNVfxt6oO3TAtuTWjGU
QB8lCZASd3ScDPjtZlQaJRuH/XhLAn6wELSyP+hp60sljN5qB2Vdi5BW4lcuslv3o9XxJ1jL5OFD
lqCW/pm4qjm1bqm52e+SxffWxOqE6NKwSbtojCAbGMZk++NKAGGUuK8o4aOf61NrkZW4fmdO+rLJ
aFWmkHsSA4DaqoPITh72cDk17AA+wxdIE0xNe6kAYiGj4/Dhnq66E4ukzPTDVgqQZwi5xHc8MLbC
+oiCrUj71RWcdhXi1+PfB5isEBSp8S7YEQuF2058rCeDCY/TpOyC3Ds7cTb2P3wYbneW/w40E3qK
d0Q3O5YckMzm+Fx7psIWEdx22l3p3jm+DZm//Wz8AtJqU9yXNGimQ7l//TyHOUPRxG06vySMAcud
gOxxOMKUtKn+tHtv3mlkmEMz25R++Lj7/fo4BfIxOidKMgoXBBdcbAJ2+ZoPcd45WapM5opkI6fK
YjUerXbklDVcZTKTyMlSkz5wSQuPXsSaQ+WmD4ZsSlBYwBKwCLrl/oLde4grDG8weqTpstKvnS5L
3Wj8FdxOvTt3yvsmvewlTUw79+0JE3sV/rfkZ9X9AGWkume1HWfcjaj/UNwOmFGwBM0TH2SyBoQz
PoZYeIJEK8RL86KxfEL6RZ+lBPytjPnDfn7+XaKJOn0Gycq/EpSksqJPdadhj7DPfiqmFYABWD7Z
OZs7M49EjjRbQQFxa30dyB5vyNMmRek8Iltn9XRovJUhYQNPSDWwqdpJAeimlMljJ8tGMrD7qyVA
EvnCDySt63G6IhAS/ZfP5pdg5H+F6TNHlxA2MauhA4MYExrubl1u9agQirVwX0C0D+rsq1N3dOA5
Zv9FQaX9vz5Q3hDc2HyOohggSj1nwcje23cNr7cRmS+R4aETFfGQk5Z7PCckVt/+t1g12l6he7Qy
k3decrIke9nfGwlC+ERAj9plUdDpeJgCOsrZzETFH5HDnLGhqTQPFS4o6RaLbtoZmvZ9sLOeq0Y2
G5G8HTm0fBF+7yQ66FKTYsCS9QZZqYoOEyBFTHgayQ0PatU3EkdTCEstVWSzH0Gu/6Na3n1BrVyf
Sh10lZVZnoBwW8Rr6l8yws5MXgnxFRNKXIdtsR8pKuQ8enU4H3QRSQTdEYu8PByaXFCKmOTnDZoT
Aoy98f256DOXpTifpmGPIyhxQIOJnM9/yZ+PrXkznnQ4SfMAorRzVjkZLRA9h6eDgvIVkiH3cDmF
9UYAyyGkss/JpS7M6aHpwRnjJSogsxwMSu4GSmGoRlVgjq+efq89s/86hYflAplOVyACEZGg2pwj
hCXqma8mdhT6CGlZkQsPT/fqVNJnTS/hbrJavlhWJFzyUbfS3CxUt1WU8tAyh+DImAKFRtiiX/kd
eOoT4VeOOLXv7GaXCMFpjJI+ndMrdEvW0IRMjD73ywRLq0xMY54JjSs03lsMJWEfNCeK32zda5lH
2Cx2XQ76utdeF6Emlg8cm2UBQdXqJniI8Bz8vZZOMzKr9hjImWIZbgh/OO/EOKnnyIBr6ylhLXQo
nQwOXUUcPV3zQadIsqCmQ4Uc2bdNwtjvy/m8ptWTdq6J8XYjIYwLAF/Yjg5uCdd8xF0eFegPRpeA
Q0U2O5nfQM9xV85f54cNN+VH1PrTcnd5j027z2I1+8QqFASfHsua58cld7FD/Ai03FSJPsryMUuI
1C9bquRPzkElaucnQSdRsDRqgmZVNDGnHZnRc7npcuahWrsmzQFNSmyDLTRhait3k24dU8MrcR5d
lvu4RP2IijFK0L5j1mPwrU/w/RBUSA+zPPJtnPat9ef0fOsaT5dlJ3yN2b0VN+RNfQd3Lrb/oIB2
D9ALWbE3zA3cwbWi2x6Tusa5VIcQvkCgHfBh/ntGkLF541nIRO+DjVGn66mWOxvBYQfkqcSrP59O
Cly49sxvoMBWWp+4f0sH91uHJTBC8KEn2zyHKJhGjv4tUFkcFdsy7/3O82Hfm6dhJz+wNC2mM42F
muuhE5vjG1F0X8SOQ7csyswAJi2If8lPbzFUNN2JyHhEaKM8p9Yul5l1P71fQOK82MVi4TmdwRgG
hTHrJGve48mykkS8pJV2NuoadSIP8KsXoKJ3lasd4ykQeqhvYdeHYmf+AoElRRX4SUsiOP0H7Uqd
orgYFwjvxiNPq+pcbtXrB4hPVlMalCOcrEf2l8JnpH8Q7ZnxaNR8FYdWJ2csa6j8Y9fe76r0ueNk
ks0sdulcewBRDa5p0QANc7/cFKgrkUoCprxpDkA+lrgUcBy9nBVOS4YdzY3KfGtzeEB6g6BU5ZXp
xwixlvo/tIPLDRnXRtoaj4LZsbGDXOlfNYtoXSTuMpP/1JdcXWEto44wUwAI8rFgJtjTrCn2z+NK
rP7MIL2ceG+bPxpfiCHAImni6ifwSVN90dR96Q7+r36YAgmvV/Ln28HmO2LhqQp6eOKy7bfGe5+d
j12vP0DlyaEwNvuV/+SCRHBjuUAlWMelDECD763mZkA6qf65zBDF814nUvXbSHGMLWBNPXaDS6Qs
dEPhSrDRrHkbfQ5t4ITcCR0RO1FbEaJvHDancuGqEr9ahkS0i0YwWAWA597FjH/Ny3tXV1ZzCTMA
uvgLhyUptySpxCgB4RwUn2PLiopfpf++PmdcLUVnfAwqt1cVUAJa1oQlRsRzIMiyyGhPgo2KYs5q
deBHw5EPOwrO+7mcDi2AwgWEVPsgWIm5A3D7GpFIDY37Z32lAajMpDd7jMK17l6n5Rx9JAv81Kaw
H/I8eXDZMsxbmgMOadqQvcyKyu1QEqDIFxWQYn45PbJvn7hKUpBPpJd3RwnHtxf0+dE2nrKsBGoB
8TnB88NSZUoEzRtObHdiSByodyAHGhf9f3+6sD/zTI657HRnZv/y91CUO3TWKcy+JDDjU74eAPpL
SgQZaqFEs3JgkWSk3Tldfaeru6MIScMZ+FF4vXXaIvW0VPoOlz/KaEPG+m8Ohe9+0+M2WN9j1btk
yX16InwNnV184aU4c2iQ4demDoOj5Dkliqz0K7KxHXoEivvUAhzQ7g8MwuIYfEZLUy9ijWI0SPn1
1NaXKJS9tlbT9bCsENw1+OAruHJ9L7vA/R2LZWPDvZFsbL/1F5lvKwdASNH/y+gqxd0YZg8GsgW2
y4rv4tNJDarwTPmdRakG5UvXhMiCOEAuOF/Ptp13H6y+lwXfcHty9JcYR4f71D+oAuWRwEC+/3xp
VPbENH9TLYfPqa9bKxQEsjm95NhkZspUl7ZTV89OiukSySCwjvHoWubA5KJD7hJkGp3+tXu+LV5z
TI0SiWCUZuFZTo9X/uKcgz+6lYcZ5ClJ5x/LKF0F2xEZ6K6J4OsatUpWnONhRpzGPwpwmqculUy4
dhMHBwT/aEu4xaJ51aB3DHvepI+LACNLZqyRZl4KfquySHgElEr0LcZoe5YguZHDreUy6cnBwD3c
OmUBWsn0gwbDo+Gxr4BcCmjvQWvQq4ZzdQahmDh7P8cPLXyacBYk1EpgtFFLpvgVzKY1M4jgsyCc
WIkdjCvUY2457VfcWOwwbK0uspRszeqUUGKeeG6krVZEZ8CDqolCvUZGkHtf6XIAtcRbwx1Aq36e
FaFB0L6bmFgkFXaGQCxhqzLAQo7/bTuisc9iJ0638uMVaVKVIZzzyoOi3MTPtOL6RzG8EL4qqzp1
Wjf0HQYvUH9ibvE1y57AgRn8OIqE3g/M8Mfg+14cMlgBuIhJDdW236ZbKCSQs7hm9rK+1XsBQyiM
MF8OwuKADVM1YJhON+l54oi1oMNR2NrAiSmM8eda37A/9AJLBM4XWbHTluCLMeyyDlnxW9h7pkr5
DrS1m+Sl+2UEvf5xN2TDeThBrd30QXLDGVWZbwKjj2+VTClu2+W6GY+ZO+fR4Z3X0Y7YNtb3E2s0
yQpBOeNfniXD0RgsOMTd7tiQ5UDduPyLWT8r+aT7b2IMHJLJbIbhx+F5qZ10a+EJ1i72QDpUR0Of
eqAlEABK+ez4FYRIJR59FBSR9LadifBDE6SWDN5k7yS2DjvW3OUxFquBVTQQScyT66qCsQSEqp4E
gyMIz01vriDNidL8CEXFsIGNRv91YMv3pbmv6btk4xzNEt9rILadkQKr3znXwkE4kCPIK8VKQXcj
ABpHDNSNqYNGlfxOGX7s9uD2O+mysy0VyG7gTDAGBbevHTMK43/I8pF+ETdVjjUArLGUQvUmbPjj
ZGx6ttT2bTNUKvM2lBhPuBPhGcxK6cxfNRVoZJ0UKHjsPSxbSdaAvlXxeVve2XdOgUJXSq+u6d0X
ySb2H9Plv4oH/jQKE4yCQMk4b0mNHMFf0YeYanO2O+q4KDPzumYGIdpPrNqoc7Yk21UhuWdXPMMf
seOCiaKn0YfKMcZGS2MOoOKh7hl5sdEcmTph3d8wvns17KXmyeLITrhaX9M+sZydh4rd76ZbqaI5
YdmMzHSph+dXK0BdcJAv473ZI8qI6G3J5sglMdRkKynnwMKr6IBnYUngATQW+x1sOs+q2Q3zAIR8
rT8g9D1tUNgF39D0jIVMGhduaqpYBisA63j0jAk+B1KvBa0KQ40LMWZzQxmp7oZilYZUnJ623E6H
IfLCBX5W4NS7/uG650GQS3wvb9l4BuF8Yic0jxxUDOlXIdPnAnyiZQT9SGvsgPmaED2/1E0NnXsq
K/HZAFxsnLgxrEuVXZJImXcdIPx+KZJgqQGITAq+bR0nJnP6H1NTVRi0Kg/36vClVPitdaSDQSAG
eL6djY/Q6Gg91X2NBGq80mJqP7vinJIyNCLd1SBEdGnL0OfYk4uGtMhXE24cspJ25nWf0JNJuyb3
uD+yuAfQnum2GZjkn/bxLvaJEJEJLh7mMUZpG7MNT/8J4Oo0vRkLtSPQTz10oAdJZYwwrdU6tv5o
ACeUczrFnTW30Q5aVwGZVsaJGpdNw/kINKS+kFGLVDQBcCWYl6i2uPyq6yOMLwHtUQgjNIlgTr5J
pUeOiMB29GPj2ec3KzDO+6JXSDHeLgI1Xgx1sGiwiBNUFtCjJogK3egu+KJxqRq3x4/WEcMneEan
Qy74VjjnBtybIbvm8RnU3Y1RpvV4q1LUP0XfV1OTRyeAkY0cYGAk6abkoniUc1xJvt4KATgEHkkA
HkIiARttfvC34RK8T3N9loQRBV/WzoU0YWeOkHUT4DUdp9ZCsDXHUtys9902IMuw1emtI0b1eO17
kmdAv+YCDCUwsMqlNKnlXHXkGpvcAxXsfklDAuN32TlU3PCdA90omYwr2VsJIZDHpFvHLl2wBjSi
xtn+LxYlbT6vn8earP58TaHZyu64nOBY3qKjxlCxCckVC/qjglkgxPRZv6pPsk4fHrO0P4jX17Ki
gSRNHj/4pn/o0rTH6SG7Wtgt6n/SNnNNNsDSmBoGnlD92w3oIfdHoyIXe4Tpj8QwoHw8Z1P0gTWZ
Vhk3bxK9C2LE97ZNfMIg0h6fLOsJiznxkqL2ct6veYBT0LHdXgm+80qvIuRMMw6cmBXaM4fulsDf
FN2rYWwDDkhxRMvA7wEJJg1r+4fE6rYE1sTPpMe26NKjOq3ETSWTP47W1mwE7F929zRo63fEsfam
UaAB4Davld903tUQ4NMiSohhkJUjji7NajAq7pdR6EnunmuFc4owBDkXY0B5kldcO/oKEMPS1F1s
l1nSUhKdj1dXM6D9roYZwrt1AEHxAzkRDCt6yZ0csplKdEFa+JiOnlNvlACp3qVSPDKK3S55UTl7
PUwy2Zwx8AXT+e4Fa/SfqtFIBrl1nlhpBIHx0V9ccxXO8D+kMBjY2FNY/G/plmQxHldkRc06/uDV
p2wxePkKaChC3VXn5Giz56r7ldo8Z+Lk3n+0e1h5qfjC3MGypLETF0PltbNxMkRnYo1lv40B3vvr
I5VOLHWeoHLwsKMa37JoRDUhcXoMiyiis2UFE+e+GNgcbsvyy3HGSlm+pyafX5lK5Vq4+/mkhuuP
rJUumTsRy7P86ZWTenqUgs3UrMif2HmM2gQZ5E/POxF8vOSPjnaq41D99fpVX7XwiOstUpNuZhd6
eRaT1gGoapQmh2OBvwPQ81Ifydaf5bIJ1UK5P688o33UquCJMMdolHh0oyVDHCkGJ23sE944VQXR
SJ+W08+Ok7qFt74zDfu2Af35rntw6KIJlWeXUB47ASnHWzfn6eZpOgeXuPczGYDEgncn5tT8vh5m
Hv+1g/UuP//B5dnuP7hZOhd5DDFOwlTp1ul8HCWqGdcIQvgHzcEoe31m540dDVCjIDEfEo6tXqly
nhXCO2I8EQDLZnZhTxb+PHR7MrL2pA/K7YDjeDS/MC+wAYi/YoGNudrdcYA6NZw2r3feVXrojln2
2JzcBdG4OmikeIfKKoiBwtQsIdgV5V9//v4O0yit4E1Bs1cW1YJVXWUOyByMrIUPvJVhDAILwUFM
7elAbDCBzyFLlg1dOa3nquQIqmDMhDZjC9quzd4pjSkVlDgCwa0WVpp7oY3StR5C1IirUnU5esCx
3lFTxL+SqC1TZUznI7almf9TyVmVVoEBO8LUHGSesF069+vHrtB/ozlvI4A1j1rshgL1UrjviFJD
OWN5yQm/J5gH9CfWz+cRXmMa2eGlhf0VZ2bPEDBozzjMUVVbMnMgBR8mPKH2oYS+PWc7TjIPQpbV
PPgbzzB4z95VfUW7XpUST13XL0Gi1fYeiXshhdc0zbM2KlgJWUwg4KMLt6Xciu8OHUsLZR9wduN4
AyyW3ija82IO0EHe/EBjp5XrhyLEG8uCrqqAKZEHla02TuUx+RRr8b6Al+rAn2pR/7bXKZzkNEQd
q06zXNFv1vFU0czETtvIYUGNe1hg7gIB86mDeHflf8j7Zn/DBEKRTW3XCVQRsqlLMsjJFn/3A/dj
3VEoQ4rIq/VX9sebCXvnhh6+KFavpMT/kHNxvTLzKCYLZLj2kQrVaacJmHnBNkRt4sT0wmlJuyIZ
Uohpi45jbVIZZcD1MXXsK1yC/dBqTBXVkYqTGEgfWp0zhcb6xoJyOAJEBb6QoftCluwYw4XrqXmu
jmCAvCCUghLHypSgwHUIf9dmeF5sjPcRRd57JLmHfOwF5rYutG3pQ5jOL3ILpyurh0cJs+B468NR
iHym9Yc9q2iNW05Tivt0AyafL/urDY0JELudkCcK5nnqbJEx2ALytqmitdU5RMmjDHk9IBe8Q3E6
l4ZMa0MdcxX7pq8/S9mswXG3g0uga2nIivNYVZ/HS17uBdb9bGkXqgfZKScuuzqbEkWCNGMjRTOA
olQn10m2OETW4X/B8QfxI0UYjk3ds1/G6EGxXsgvN28Hhs/siWMLDFIPZqc4UBz6V18nQlRVkPVp
YMO2hogMksP6cx4Ogi90pr6++0pxgMYe6pH67ssRDtJOcGepmVGresVwokM44HSJRzKwee45UJwH
lXkxYlIx+sS/2PalZdRKc6LK/kvS6QrC+F1DSDJNU3Z/hPE4bY7wZvTa50wZFycVdqKW4ojCcFsj
rxu381mH4HALYvs05tmpzuy5yhpxe9vsKZ5mfO1Vzu2t8sgvqvccMbW/POsg1PbdTdamew0TSGGe
QDzpLZQVqkb2Jnb7czC7br6f8lw6ph4rthoE9vUKDPiqVSPgpOE8kxcIlihpnnkdTevBjUFVdKFR
nnR0CEi9/g/U2OdSf+ZC8FjYLfLEqveubGD+P+z1rXTunvfxvh1ht44gNTzgOaTO9gEGh5RMx5zz
DymYPu6MkyP80tIue1CwZsxm1YPVp4C2EyswLnyrCCW+5jduPGqvUQf35t+/9RGcZup/YpwQQnUF
pnogr18ufSmNFv5TQJbhFmU4+2bsxq8+VNn8t3ORWbWrnQoEbiDkqJCqmr1wNCKQGm6HetvmNchx
lk6eSYKk76/Zi99/16vI+f0w6LlZ4P7LpxX3cGeFmf6s5eOJKtXafp8VZPZiDW3tjtBP6p77LfmW
AlxN+rFo/4G3HMusEqZooWwGvAUWMJW7V2faT84EuoyMsb+RmqYiFhjWVmWHnBbVybQ2ZuNPL9qs
6Y4dBx393M6cj1U5e7Xo/D6cudViHSrDx2AJVfrvsPOqvqJZ688wBKOYKy0kdbqQpqjSG4tbk1dW
U1RSfvEDabgPv5FR+uT8WYAR31+J916YsVn9vRUzePd6dDXgnk6I2TLZFPEvbbrtNEdB4d8jfU2x
S+LceyMb8+6C2nOuj4H4J5WG+WUgq9kSSGbq+7sHsaKTIBewCOCQxO4CloxMod/ofrcchqvTgdFC
SYPfIq6/PrPOG/gmqhLCvH72mX4D9cR81esz7zWJMBaS+AGBWE1wcm7YbUW5JQ6U1OmSY1uCRuH1
ppTQ96F3y6CFr3EFMQvLR0djlf5uLZgLewSDurGnzdWyV9Tgjk+FbbPcDypxkCj1uGKnvBpkOSRs
S+uO5Q2JGOS9lRt33xgRAxZvr6D+kkfflgfw9SztYNFV0/hxEyi6KNn4+R0EUkiMKnOqYztXIfFo
mHthA/+VwJ7dbSetewsgwQcZzYpUHUzdr00M77yyxsplGqN44LOwdKpGqAkWxSgrlKf8LrgJtec7
W8W0yoazBETpLFRdwC4GQULREFz+kbBjG/O5sUHV7E+a77GT3iZyYLx9BOXwUCl8cqDvt2ZpxbS+
wckb+3ZnwPC8f+kret2xmznyIIM0jo/g5RP3FnIZ7ZVsYdhSQt8KENc4BdlF00WLYa7Zmj5sKVIC
FOihgXtNYcGk2dGCREIzi+O4lyqmop9HyRv7Sth3Gg8CXjPpD35sH3CWBu4zPqGePwkkqwR7E3tX
ecy36Uf6rlM90OY8c62ELxSu0N8tePNkGnsXQwGmHO9+Exnb2htQ7aqaZ0o5SCuX6c4Zn1vnflsi
HLUfm0ur3akAwfqOxHwn7iz8eNymdZORWYwDtYI2bVhtOX4RBDI69jfw0nJtoq9qHgyn2FjPOMVX
NF98EmreWYR/5/UGnlDeixyRiTzq0Ym/1+z14UtXwHRfuOE1SVH3VN0GE60Q7TJ3om1qOuNlz4vK
pZ76pXxN9lAlsJHbjVsgW/hjxqtYbd8QIHD49TYvgYfC8CsmXjkPqom2y1+DDYigW3y+diaXTCar
HgB91QLZyfQjNI3v+1gPLsC3FhBRG2DXaaNrfzIwQKtGezE594iyp/3uXywm/pwTfVf0jt+7hkEq
1kePcX7jIkVKaSuNLtB2YFAEXUKTQzlCu8spDEr6jzIHyQacNuU1rd2owfR9etvMRlCLaKa//NrT
FgFFxfS64Jfh6HYADXNOsijc95gN3YcUsaBo0m1M2cKEN3VpVuj1HMMSjBKCGeHeXIKx6oLyo+rb
0ay1c2qCnb/ykTGIB5eapCOaymM2zzWLpMmjMR/D4HkasEQFlhB0nBguZUKgH9PdYvVg+1aoTKo0
Sp4efLogo3w3yabe2DMRl9ZcJrFOqapsJ+qBoIkxf0I1i1uxcis1ndTrIGWhWGicA3I5+NfNAR/d
bJyO2P7wWhTWaj9sGYM/f54H7/IMrn/gyRWg7LaXg88hLxliFC3c+jUC4Mw+EzWn+xQTatOOXpoI
F/1gbzGh+AmO/p9HMJUxfZ0BDiQLG1iI0ezVgzIHbRd1A8uNLu9WZ3yOvYzw98qi83s5wJo74qn0
TsTkC9RkLMRQaaFQLRBgtEzugAqNWmNMQXw8Y72561Wuu15MMgD5Wg3SkdkHDaNeFeeUeaVVKcaN
Mf63pMjLo+r0jcsAfhz14m+j2OgCHP9UecumkqWpm0Mw522fq2E+1glYHd3uMvcL1hwiSgYchaTA
FGCZvUqY3FyANUdheBu1Eb8xKxqA8RuHFYr05RT4vLw3D7vNqqOMwYBE26niDe6+hJKHZTeNctWy
MWvh4FSk7cU9Slx8LjpQHupOkpJ77TeTogZWNs8JGUnwLwW5a1ALKEr+/Tmxk2YAemgpzf/Bcqiu
zQ48RYgSMGqGnuBYeIu9FjKFqePGgxRSUkZrJiM4SLfi4rKZcJ1VVjgU7y2AL4t2klKG4ElXppci
+sLgXbb57s84CHqiIhNG0TIFdEMWJp2cYIE72TF+GaTOjJl35jQReNYhBP6G5A0N1VJd64bQ0QQw
e1UDGbRbvwnGG95bpC0DK8I+jq129MYq1d6ouTekjO/S8QuJTDtCxArq4+fF3pLoZwfjHuH6kZfG
JHm+q4yMmvPz8zwdH6/YW3AczMqvw8h3rJqey4a33f1/LXo3mYrUvwBVWoINFqNQgUdekZpK/jdF
UZPLgHzZCtoxKNOZ4g==
`pragma protect end_protected
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="default"
`pragma protect author_info="default"
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
ga7z3iGMhGhga7TzPGleypVOHJn9S7KEP16RJ6j/y4QGRddc7/SJdXJ2zPvm8FTCqWlJhu6/s34X
gPP3kw7dN1YdiZ3wZ0Vzt8uhC/B62KTkMGylsJT3Hm/4AVsby+VuOus10FHgOgp78G6FqJDW2hD4
FEF7AvpJ8kF9S1ZR/yBaB9R5/vEzgMTG6H0b1hzTpBGPyaW1S33KG60mDs4uY1wSc9WkIOuDsX13
gE5v3E3AdV0s35W8mk90srPFan8A4v9WhQvKv0pRdTPwajKYNoHYw9l0a0ijfdCCo0SwbSJr+KOr
7KJQNnQdeGn2Y8dg3BGFPO1H0k02bZuSqUQ8rQ==

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="GoWin"
`pragma protect key_keyname="GoWin2016"
`pragma protect key_method="rsa"
`pragma protect key_block
dBwrqXpaPIvc4b2fzIcAYNKycDBKm/hw0N9OirP+O5J0w47WHpIJLrz+YZdtlXZ+W2OT1CCdKga8
l9q6LpHNXfMJe0tSBaUQJS9kx12QCBYd7pz6Zz4XteULmwejqAW/r/1SNtjKdsFfgoOhPbvsYv0n
RR9WE79+rnvNSo03sWloLz3If8EsTQUj+4AuHA6W5eeLCFFrjEJDELred9ftNf+GjbKQ4DD9VT1l
GYpqKI157tMW7VzaYctB1tIYsZm6N1scQY5/pen6aJE9XG/GVJc/lUhiKfjKkAB4R0V1b6xO6o/L
Z0CvpttfY2ekIVc0VuCKq5gMTfn8BkW7RjZNRA==

`pragma protect data_keyowner="default-ip-vendor"
`pragma protect data_keyname="default-ip-key"
`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=9072)
`pragma protect data_block
3MLlIGXYAu+SNVZUrN9axPWxB76fSavWP25CyQigoZQ3T579rH2tX4mOroKAFnY6MCrE4zy5SoFT
o9pFhWobhy1JNncmCcy/a0fRL9ZlIyjwjHAt323ZL0R5G1zw5cvTmFWPoZX0yo775l85Oj07XBYY
i+0FcCRCKdgsQGwhMUnpc6ET4ttBmjQUuxB6g1Afy5ISJRNYs77D5E8aOFrmzUzDFsE9BGcX8wUT
bT4zFmjkBZBQ+KrbdhaUiVbninMVuzKJe0egFOCGcc6CdMPwZP2SxWGkscRsjPCAUdXGIydg5Z31
50m/zUoKITRK4jViYvnHt4f6sELIUTWEwPvxSg4M+j+wpDH8hMQC98bpm495w9Lz7AbFBmLBe5IG
17+sbfU7k0MY2fUrDvsniZvkyXNkbKvNrkm2E9MAmf3uKtqsnMU/tF2um9tYyMuoXrnv+cf1WHME
rcGa/NDEnGr3zL8P+jWgeThli88TgswwgsRldtZSZHdEDO1R1Eb97kPR2KAaazYlo2Q2STr+5F6V
SY1q0ie4TtY/nmeVptSZJNGauW3hhgmAK4fuCh0LfgbkBsnHNuCX8t9sRAwVUkoEOlvg+hIeL3ch
IbMuCTBsi9ym1EZ2NwdIt6YMzhAa6xgt6mL0uQSzppyrK9CSimYyzPbah+kviBaNcZ+XJClYLFwg
Dt034rBFaffea3MI9/T6EckVHZwmBgwvpnfxe5dIdxVZcMCrn14d+8gHoeJtodrk7RCejHv+C9Jn
yRjIaiu6w3mbAeAL4r66PbCB+S92jMdnwdBtSBcwI+pRfl8Y1ZjnMUax1D4+e4G/2vS04zWOHJPK
TAm5M/l7TRLujzCl4M5tq+MN/Sl/TrmT6Z4/ZBXtoFpOHicvprtU+bB6bA/TDiQ+wyauUCUWMDnD
F2sWssLTcUSqWyGH8nZQJkJU1GRznsjpDp4OUZFEoGr1SIfqUXOeUdRWE7kTsTGtuLLkFRULD9ZC
icKwOzgQXLWvy1haIHsyX6SZ+d2z16A+qjc4h9yGuTAjU8NLa0V/nk/gnsMB1qd073hph6QLxLJK
r4sFXdYNYgCk5RaS44kcalofpqStJQULijgevhq0IIAiHku9ZgDSCzWAw3Mr5M2bNizLX2XXA2zw
yD5SKKgh8NLJ62Z1MJq1d/+XEurLezROXf2MzGpmtx5eT+YNTMToyw4wlcI7tOteLNTVwpN45tUQ
B+wyQRROLfJbya1slSCz3CBx0TkfIQfh2iiO78hl2uIlnw7hygM5cDhSSbRATA0xa7ahqhvOPN7M
cHlx2JtFdxdsqSaZD9QoJ639DDyU3Hou+ECwMn0csUSwgAS8rtGVdP0Of14CplgwrGPXstO6akKA
3u+imfQ/w8L/PLKXBmZ4JDbURy7k1H6RKbw37csxd/ZvrS/pSmIkcNCzp/c2DuOoQ7gmrvF/T6P6
o66nwV4BSbtkXVm1Gd6pj8kuzFas4d8qUgIJYtO74n7f/EHBC4KRyKr547xiGiwhk9b9qd0mjPKY
rhYsYy9gXuZh3r68RGneNEq01MvW6g9QFwK1ZOIvZDYOR4QWzSf3jaria7TfeR04B0hTDmN2pnIe
G0GNQyny7szBaDLk+3oC5dKi2x7IBMiFePNumBGpRQwF3BZOBafJAtsThr6J0+IuaIyGTu6q0CRE
pK6/stbZUIyDHLZTtsEiDvCUoqJt1Nwycg1jZabyqczbNym1H0NA+utNZBXESxVE+E0tL5xp64UF
6UUd+qxyLwKovERkzivDR8GuW1zTirEOV5S4VxepjAekJHQRl/DLLebsO05p1WmBlr64t8l3I2Z4
eBoTyoAckywhyY3Hef2UK2jwBO8dnRLD1Fu46o95g5M70RM/CdS1OdLKSF5ccJEDtzouHFkJV1Uj
jF3ui454vNAg2ROOQ3kKuyo5BsEY2EVCu3TpZq4c/q9GQLsRGPOnx3VcTR+6BZb9QBmDwr5qk+/F
Mfy0nKqqzp3OK73AWybRMjmJczTm6ffP4zxEkfUdzR127EO+OljvRItBn8LSuKgqUpIu2NxDCg+f
A8xmKgcdP5Vj8cz+tus1NipaLcnS3rd6rslS/DaabQM/fOpx4ERbftZUSiDhPxRfGlVjhYH1zMEk
pr486KmY6LfVGaqc2pCdgIkuSoohsNiPN8xmmK5O9HjxRm7IYdaUIvotow0YeYsJys+80/gJB5s6
cE/ss5YkBWNMAqtri10qAqP/lHRchjbTFTFInn1auRmyFcN5WTjU9MqXhbmBIpJrVs6hQ8bjrGbe
udyynSp5mkE0eE/e2v5I1wi1YhxlXU/wpSQkq7AW/DgOKirxvaKomORblPuNuqND5ETjQo+jpEPM
80/aOZIyPqN0aWmrTJE0jsjxS1AJ4MOENCzTG523Wq1bgye8XzrN4fo53VpdHD6EPKSh7ZgGV7sq
giQ8mzKHA5CetG2XXI6zrPk7Oe4z8m90oe+OF3HP34C4sTOp/x3Y+GqefIC7NoHPNtvs6PK4n21W
QJDfypWh5VF59VtNEgflzAT2wYDVtih7VEgDNBwrj5ychDhaeRx4+0dTJ9BZTa/Q0qZqOY4erpsq
jvneKxGNPh7zRngog7RWOBuH1Hi9ahuIiY+gEC8RxoTw0q9WCloHfF6cK42Bey41W7Nkg8Ic3W6O
AV81HlRcI218/r7yKU/7urKe8KAq0lmfWI0uIobow6NRr57vlBBhnMIl/DXynMAD0MicHsH1Dhyn
h+XWBoQuDUWkaHIh4zZ/+1qRMEs0NnSiSUJpOxoccGc+tyhoKIypXhHvUevk4IqtTmdXqAG9BJVV
k5OY9fhhlE2OW/ibdkZv1N8TAqzbACTxaJsG4yd9IXNrWQH3memdIJYipNklf5EjC/KvbTm5tyl+
BLxlplNCoR4T5q2klsjPNTl8nKAiMYCZJ29rISm9ghJjvtpxxC7iQxNuwy8DpjfL8Uf4MMBxii/H
GSJtEZy1R7DGqeOvCIAWAjS1+kkxdMrlh0x3ruEo2+mWagYuF7zcRwv3TrcxsdpZpxjAK3KuJQ5d
X94lkof9p94Q9FjBqgLyhEjFTPbeSIdMHrEiuPoqCq/SHstw6UAe/HyD6+3m2O2WR1U2m9uPatvm
sJxRvmVVaHWurvpn1JNRY5/mpZqXlkjzuf/rk4eL7YaveH1F0WX+Ql3Pd0MA4RpPOCPoYJ6ooi3X
oVoBCaBgNLwuE9nJoaTWldtbdFa4ZaDZk7rQMlAKVWXu5XPEChTjxfzXr9iZw8Qdf1rTNBPLxMWO
LS48BLsmr5GXjy67UEUXHgGbVRrUX2AYtWS9hX1O9CEOcvgQiFyWG7+HS9TBB6SQ2461BLLzDSIm
tHQ82QNlJVtLqGTo0WcNrWtZBNk8qWHaU3vXA5QOlhzZmHw9E/y6jLn511lV/OUgJnhM+VkJUv5u
1GWSh+SGQ7IGzBlp1mAMXXSKsY9cSzVqiU7ytCkCfz7j3DJH5ntdAicnI7krHr+QdHoHVl3cPRNN
NTik7Oj2TIhkPWTVsDBGPqiRUwIeX6/EI9jZpwpEEOFrirGLMXLQlE4bDVag+ARha7L0G1Qn/UwS
ejMGqfZQRAgKydtDRMPe5ZVBcXjxlbFRxDPhda1EEu9YwjoxssFUFYaTKNMkzgd/ILMYuoWISXaK
+L64nS9GUjgI6nDexUaG+DxiNSa9V3et6jDkOQxxrgWcmQBpkk37KtycdmM0jrStFP5wmOsnlJFp
SCGPeuT7Jqp7MdnYaR5o3vKVglmGTbwjVEyEhlWMC2Bbyue7NnT/dyA0LgjQbOF69e2BR2bdmIIP
aBoT0VEoRqavKJW4VVJaM54H1gcMOvTiiwzgnJDFqLa7/UA/7wMiCGu4uBnB3/kQzacm2hlKuJQf
T0+vWNMiVBUy2cr3ft0/kuEG36VBq+hWxfKK49u9O1qhxvIIn1z1ZWZZD3MHuAZXojeGQbtv3kru
U3XT+pJVLh5oW7JXXxSWdaz2//oEhs7UgNjE6GxBsIMlGPBbkJ/ycx5yfyxee/gm59BlN6y3qJxe
INbnePJ8joraeLI54HYhmuIWx90XFHYoDJPGQspHtIFbLkbuwDmzVGbD7LA5GRjFnNUrTZfAP1EV
adRX/fDuSPpw1emPPqmQZH5VK30d64GZveWzK9i1yfrdv5e65TEzX6LlxttTYQKkEP+dtczwig//
R1YueNMWN0TwjToe2drBo7oIH3dvjjmCJGzj7L0KVXsa9T9OWhDmY3bFcKwLDrLfrOm4R/IuFEHK
WOdLDSei1hDzy7wy/K8jki8xgNIqCnChyI0UL0h7MGpoJZmBKzpmB21NrbYCdS+XnclyZ4pPkj97
Ylxo6BmW16US+sj65NAvt7uBNJHj+3T8wr3qBqSrSQsvZLNHSB5/u+5ZrPQSNqbhhjQv0NxUm8rW
8mlir3nvxXFJPZ3K+S6GI2Qwnf2OY2Rw6oMPtCsWx/sQiTfPQtb0pb9mnbOcVNeiEbHXgFZ0MLGz
HSxuKW1kexbxYUG3eu6vL1dlUHRKIQ/2irLYTwymVewOAwSODl+75/uB8Wo0kVVvpXGw/mTINAYu
7qVxHRYXpj/ksW4pfMUjP/9kM80OPdcSc/1g9yUPA2RX7QkGwH4JCwwFsIgv1mvu601jFz0O9Bkl
0PpkocFdGAcJZC9DhmjGWZD2cCN9j8QnvkQzeLUERyt2rqFfavwGkaLpxkfrv6OpLM+hpop9o/W7
f/p/JrT5qiANXTGmqz3ylmPoU7Tu4TIZURP/95dqi3BHf6QvnUPTKGAl4uafN0PLzeEkjspNN5/C
vni04/K/QKDpgxa85gtsasDqyIKmwUwKZM9db8gdA4mIUc8FLdgw9dfgKKI4tgB5EpPMO/Tj4lis
tqjm7rIoMX1dCl02nm+cc00Ed2SnpCSRajJwqkmgz9Uw6BQK5BquKLHcV+uKhZLq96f6F7NxXbnC
VSmpjLjMAEWoUhzZfYGWzNZOcaJaQoYR9IXGrPsoNr30J2p3o8wNrqGikw9KYNxK2WvLCY9Mm7xZ
ANoDsp+v7SBkr8eLvaW46it+Y7rYG5klsRcSUw2nGHzcpwmn6qcJp532CjFhZ8hmxQdCEJZIwILp
uVzRdxU2t90fe9mLoXkrhCopSuvSplsAbKZ6yaOhsSOu4PuU5VUVh/u6OF/PfBHMdXgwxU8FGb0y
hUR83gXciXE6dREXeQKuXfCaGYRt3sEnSdXhFFTMqzCvmb7EX97OWDNl2ogFkF1eh8vEFp0cO/9x
ayCzUdCED5U4SZwamqb/MDo9zUz0PLFfyfocYTFS3vlN2VJ3g9+6zxksTm1dsSso6oHVH8ZJP6wd
KIr9m8QKTd0FXZnWiH8hJg6E73Ssrjj1b7gwI40w3m+jM0O4LqBgHZctjoM+4eYsfe85yhVIUyKV
Urgl0O4NuR1uZsW1VMGVtyngNkI31gbHIWv572fxN4ikoANmSxhGNAG8/qCWyXdQfJUNELlRqqQa
kAwhWwDVJZ+k50DJZTz8jARz55BNIjVR8ErTF/GuvisBZVjiueUM3GW1QUQeP/jr86MB0LIYNccP
7DHwyT47vp2fhU7IuvD8FiP6/DegR7eAvpv3T+B+xcT/I0uB2x8fDgPJw1/b7F5HfvZCIbNb5SVH
Tw7kBYyOuTrwFrANCDbsV1429WaRXUdBnqS4UbNEGIFXNSPuHpR13Ge402Mxb5MyuIoWP6pRx+Eg
Pj+pw3+oMLd+I+j8zxN+qdK0FuoI6nIHh8NDD61SHNGXSOeWuJ2wEGqziBE6o/rm7lnw/bQdqxSR
YV5Byzql8lSKdW32uiMMYz5nKDMtqxStIVSJkUCxjUlJ0mnGjcnXo5P7leZKY58LPiS94oXhcC1O
kzKxrKVJznqpGM6Eln8v0BX2ilCKY/b4oLhLU3B0u+qFUU2olYnVfQhZM3E1Tp5gS54P2pdf1v7c
KMuRwNntpy+X5hZYMgazx7Dov2KLO0FXoYNaiIj/o15wKmxexJw2MwilFA9cGzvh4CMHx38XNzKc
wbmBHeWpHQ2ARcOylDwPaiSrZ5E5d47fg7raWfP4ysjybfrEWn85I6dCXk6w0qhPvAXOiW4AZ3bh
xgXiJsP7o766J5nn7rYPh42eWEfuBRnR8dh4lgEAHrSM0gB69R5KiLHVQ5/R4XG1QSCw4SsV5Wuo
ths/6EB8J3AY3AfdjIkHCCeVbt5x8c4K68sXKhTR+ifR5K+G5ToxIAY+OhoJ54flErjCOsmF/Wiu
rfX2Wa8sXm4npR8kPiC5at4zYcE4qRzc0xiEcXBo9v8uBV1Vifu6gh4z5HlYIFA5dGnrDkzIlSIK
dYpVB9FND7PXET8E0tDhT3Flaubox2Hq5oXdATN8WCNhrjM4V/hELCobdz326sZQhR5GUkDcApny
8Tu4F2YAlvhn2A8Ni4Rj3USuxSiyNiEg1PAK3+1XmtcJjKSIl4wJRNu3+Jr2xP+LlOpkl124rb6J
Je/Gg5bnxJndk1c/DuCX3w7v8cZrwLv1uAZ/6bzHmHGswjZVzzR1xNmjDtRzChlCNkuAEz2kRbLx
TGi4H0rYWZ6AR8ZksqJiY4ufxrQg6Ldr8WBUJmMvtPmytfptUDr2j2sHyxEQFfzzya/rhjL11VKL
N7QNG5cVC5N31XO+mpdD6mn8gvddDzOl/qRc6SuOJsMjfPTbzBexpAWrLA9YSaGy/2R7d9hDZvWH
f5qEB1TRWgjyyKuu3LEVeIMTJgnHmeCOujSjgPByFLXLpFVmjFDrB5Aq8cu3WtWI/NfA7Qem5gy2
xsEwm5qpaMi/nT+K4rQPJ1N4gMikPiIoIGI1I9NSxhJrh3PeUJNOh4qrXWU1Wu/XMKwZnPCe9pak
HvHKNuIrD/jHS7WIas9/1iLRBIonDsenldC2bBC28pf5z3WzOe0WPpYYaGQ827RaH73ls9i955f7
qkA82W14/tV1nEVK5kYtL2JaPDbUU6Mfq7liEafhvOXdTnHAKAykh9k7HNAniy5DUH0nnOe3lVjG
yr29Ha3farSkRstToaPVDiM+kHJ8N+TCwK72uI7LbeS2+2LQRlVmYo4X8PY/ASciygc1olGkqFh/
qMNFN6cO7zZhDXiCSeSPwyvjeZXiiGBoH4a2w8IBU2AX7tG5MDMkudV+spTesytgJcAiQs6CpfwF
XsaGajW8R6h291d3smw/AY5JVSjZsYTSvsjofb2Zxm5nd5iL3iWJXoeWWi+3mZQGkXW2BMHF2CVS
71igJE+ptLEY45GJad81yapgU4axkimT3BMSoPqNfhxO5OV3Ta3odZgdYhdqnP+teV2RG/M2Hd/H
E288O8tfTHu90FcsNy/SgvOzLmoPcd0/jHLd56BDI4zowvJ69W1PZyNi2AgFDDHSY64wVDAD0Cnc
6nomSA019TnER/cjplfR/my3/bQV5gcWPTh84/J5wculwphZJOuhElTGmOEhV1jeyaq1Fd1hzTTs
lDb6D1sOMQmeA+lhr8nVt4CThr6LEBDzR0DwrW6HQCfElBCaWqCbnWiKiR4gJSIGEzIn1YHKLcCu
LfEe57KAA1/tUdDDJawHF9BsHlIPOdLTLTORxyTMSOspPtX9NVSGGUWnVvU8FmTNgyVplcWAXUIT
ee9Yg1GI27KLGOkDIezcY4sXmfonRF7zo82INxyaGwCGcRsv8J0VnEuBiejsOBoyo/8OrBH107B+
4mAc3+SyCipuEv1GGPGUbQSbUFhd8bAFZSgTVO223XsnTnv5ewREPpjR9QrBsdWdEKtHRSxfwqbM
mtPlrN3vUor4eQP8Db4NpsWWkzKRD0rVDSpXhpK9d7HGXIHpk4SXGSM9nTh2+e8N/SFKI9vr5mx8
NwwnSy4d0+wgkNtmxRUXUa3IiPFHU/+hE3CDn/4ntwb2GlKBRD6Ae6Y1ehUydDMTz38WN6cs7mwv
juVogt75j5Nk8CmgaQMwbkVFALve36moW/zZokz4L7mitltlw0/FYgtIAe3hqBryx2rQvWDf0C2W
Oh4lru29HTO/+aYwUubowRlHDa0/8At1XdjjdkOuy8rdPtGqpI0CZAJ7/DqNlAPa0gSfKT5Au7kP
YjYpg+Od05YDKTRHtEL8KTagsyy1mcf6P7W+75CEdG4k99e3J2UIXN59F75xz37cnfNt2zwWo8zU
slA09I2lTSE/zMRFXLwpUL2OZTCm8sTOfJaF59d767021lvzPdEnJkGrV2e0U4rQht4rm6Nx7NfE
Ki7tT5Rhe7FyvdRAxRhjmY1/2771QDsWk5mnuOrc4cZz63aJ/cxz1d4UJNa7TDqO2Zinpr3SbAyb
6HYsI3502PxmvK5mWOxRhmbtA5dcuDOFHSCvJkJn1Fim185yR3CbSqJ9mnavtlCY+W+hHZSUVg8P
syLhpJ0i/j2nTpJ39m3cYrFYGqRiBRf3ZDHOn3VFxfWqXpo8WCpeh2cm2yAL6Q6FBMulgN5Z9gAt
oEvw9gP+CTbAiLK4q84JfvUWssnxx49+USxDBjb0IlqWNFGpzv/JQE1jhgELytU0IsPHKFXXug8G
TXYg8h/HyNAKbpnhDyWmCJTS3Z5AfwHCFT2u0sAhLQaeDVFw2DU+IHWOcnkSfnbHElFir4Hfu7rd
EwOcYOgMs5rDiaiTrZwFkK3CKX/1kyMs3S9IgPKgrsXz4uIHvTMzZ3hQYXTC5Y4H9cvlN2Ax/ZRC
0W85mvpe26738kQ52yzmvf7eqJlgl1cNSNii+RWbbZPbk3VhTri/nlMmnwYMbD5gjWBY33A5gqfO
sBDn+F2O6Q6rk4M5WBHKAFleJJdf5IKSkd59TUsiDZvr1UFZCv9Ppxt9L6ZMPy9644PmqeX5TVzT
YeOGylwSDlWtAImiUHOWL3hxFR3XPBou7REWQHnXkRURf+MCBbhOauPVdHfwNkry3/ByP5JBD3RO
0BbSaWAc1Duqhmfy6me5oniY/6iQg/rrtyJ3ZG3U3qLgExk7tn+qxHRVV7sb84TCUojRsjdo+DSN
gk0uEfGVS320FuP78CH98RhDObVqWkjsjb8HxVbFShRf0wHoXjGIYPvSnKrT9VhN+VQkKCmUF7vP
48eq2mtrbmbOlfdkVMSDgUjuMHKhpN7/X3gKEQRaB8ai+luUtEXTKgF6vvt82XMOTswnQmanMgha
0ENrZ28dHSwgE0Snob5mYlafk1QsBazL9KuWopmgb4WsXVR9HxAkysmOa6QShVfpMXgF/lurt2eK
7zG9GMPp+451cr6BwWxmWtN9F30ZuNN26EV6onk+WCuwniVYsXJu5GJl2eATWA7gT6yNcwlnAW3V
N6qJ5Ce802YxQyYHGqr/Dv9TRswto7rNGkIkpVTE1D4mO7zyr4Vby1s/0806/bme07JVbOUotqbC
SVbJ0/W9m8tcKHd8jguDPJ3Wo2Irur819WuhbS9i1LjzNjsckztEWJKcRuCslVYfcrM8VIH/r43M
WxzbhyP+bCshRy7wEImhKIWowgsqM2NUPjzM5GY9NkDtf36bZmYZjvqyA4iXuAy+I5eQKVykV3GV
nd8rbTqJMumcSCIoB8T4EiRkEdX5b9xSrpBVOHyMv+LYnk59mP+7w8WSeDfjkIGuUPpg115vexWa
3mP3L8c/qh/AAL+/IT48uiO8fyheRJ2IXCSQwe1KgTibe6qeCPLnPWg9OutX7ZOENh3f3C9HOPwc
G/Vdf546gc0Ao4Xg9HiXlbk68HCRbcV8SrazEXi3nomQsiTxjv3ZDOQT3yZREypy3t2lJp39xG5e
x9kMEc5NSczN3Sy11zER1sNG4HxEdMYATQaYUaVp7gctY7aRUFeQLWoWulNSVvS7+GZOeHMkHw5/
yRlZwGc+cbBTXZpE+k88139MNA8KTFjmInQ/pSK4gRsUKnOSChFGfMyVoxV3Z3603dBO+eTDGCIg
sqkfNZAlKZy4ewZ3IDFw1R0HQfctegwFKqK5k+b7qfP8TbB9CPlk2XYNoaQ4PV6fKlUOZY6lDZYZ
DaNuEsxmvI792YipnSqZ+NyjfOyyCpH5DXj09Ol1XKNESmxOzpsXSaHKJxV6Dz50wZl78nfMA4WV
uJnsePvE1g/OGZaDFZX7pPEFBcHzHoQ7wa/lPUlxhTuDYaCkytVl19ZJb74X4yCD5SCY7eLuOZ5J
f0zj7uwPjnLMu402QSr7htXY78j0+MhoC7zi5vUVBeqeXvw7vmsp0zxaghJ+DGJEFei2+ROSKqSy
yWvn3lU+b2GvYmpnTWY6XB2MAHuAriIgJ4ruPQM7vf9Xvmc/GolxsRVr/t6UH4tl+67q5X+Qsr5e
eLBG4eWagKTrZYhLeeIhbsYG1ZuiOGJYVIub4e+StYBVEGtCfLzB/fJAsRESKF982kcbeg0M83t8
3UYhH3o3OE2vQX9ez+NRvo5IQF+wivGT0SK55QeQd/fRktmwSBHxIiB1hQiWy+GPj7hwHJs/SROW
8Ul042DLYuUKLkfgKNnWp6A2QkPGvgTaZI5mD4sU6okw8hErv3KCMrtT/DTepa0vSCzaZkfz1D0n
0/6wdQ0UNam4BKxH2AC8FPyVcbOdzlZNiNLUGjDMMIqoqDAJqK0y4gykOMgBn80S97VestIWSCsn
AFFReSu4bCLu3XlH40qljY6wbCw82dEgX8zInQ285Xyr9H9BnpfC0yYVkuNTu5a8qFNVEpc2FW5N
1xHep8yYN3nWEpc2EKdOzDiKYpOzXlsmrqDY4lgGiQHKvHzYSMzlBUgQzrr/eaKeeBcg7lTkXIS0
uE9xM1Dnxrjz4/NooqxChQyRsqNGIxGnTDEZkkNesW5drt32z6ILExYiTPVzNAMKMkWPxLrz5OZO
/RDWzzMteLKyzGbRrbL0UTJqJ7KzUIFO287TnxLWQhnmk50OZ1mk/ZPWebYjtORDeQ/ksyoAcsT9
FOeAx0Wg/WUpMjUC5rlx+9nQYQ2rVVQ3tPe9GnH/AGm/SFUDvpWQ8MYFua67HgTCbEzWJM9796Yg
xff1U8MwYyGKMajYwTqJCx0LvDlAZtH/s4Bjab0Gb/aRN1kF4mE3tO24yRC0DtRyGX9DV7sx9T5b
5EghNagRvM0iftiYTaeJDEKZ95sx4pV1/ITAzm1qeoZad1ybAiiGeqmAzgDuciavuVP7TtuMYiGj
DqxdbI1ay1UVo/e4DfY1Y4+uu/EtFj9DLXKD1jeEtkYPgzgKIW66JJarx/6BLgZX6ES5CkvhU7ja
B3FWagRY5+/iYjRPL/R47vQq/g33VIn6pTp78y6Ez/uUv+LDfGe1J6TuSdZuvhNgyeU15VnRKIym
Lhnm3qtqfv/angAozu26sbPXYzWb38h4dvZGwUZVD/a23013aRTClLJy+QDiRaxeGgF9bnXh8jfg
RnCAYeW0qRvv2DgVRWKFjUGkJQqRfO+wMd+s+iY38Us+wcTD4qWcdW+SgY+7gvA9R60FA9g2Z1MF
c0XSHj2NKu5vr9ztETZjqGJ46nkpduHBoPL95u7CaHDfeASF6yoWxgLbDswJkfLuPAl96TfeSMFL
8VG+f0VSV1EN/CL92AQqm0n6KczWCu/SLY/8PmY5sOTJMVz0dvRyV+gZBbRSPtixs6eklHCOMSzz
pekeY9VydYZEqQ11cmKULGF5/zNgA51lHjU6rRWOoxTRtveEyLiPz9F9zOfSJElhHH6b1R+MNkX4
WnLs82rY/3I/rY1nTNvTZcvmqGURL1GdHLE/c2WwSmWysp6hoitzNoi9stuE+6IXnuDahIvI/Paj
AjxhUbZ5TxlFZ6RTbaAaE8wn7jrp8wlBb9KVfw8SliiEYExYhdbC7X3zIr4+pR7ZDfxA/sbWx2qg
IjSSJkCcjuhnvzdLHBaQJrN1HmNUHYSQUBL6eolvzAzISiAdRNbDdJEtrYD5xUysTi1SMvSylURB
gWywb9XtPlZMnqMPDgNLpS8iL5zbB/mHbQ8HnYPXgHd2d8ecCLMKVuyR3wrU+sheD6NsAM9E1uL+
w86Z2P1C/UZygh3aAzBFK9/UHMAzM5K1LXxk+Gebn4AyFohrdVamFp/cljywjlrpVqFC+e864pGs
fuC1ghoEq7pMFhUOiiLDLI7tmw91bX51OD9hnarCl2zJmpjwLQ4dIKkexZFNTilP7hI7dw3HxvpS
CmVns1GH6E+t
`pragma protect end_protected
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="default"
`pragma protect author_info="default"
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
FF92Y2BScS1tYCbOJ6nl/yrS9tO5nLdkcinIUmduQUlX/rEFHoa3Ivyk0aB+kXloe21LQE4kGkQ6
Q9+cOvbtZsLXojH8eCz5LSxZZmj1OY0HgImQvBdW/AXKvPSh/8qp2AkQS6z06aDmakr4JM27sgw4
e8FcV4tuRcqkGs7bb5nTeggXj+gCM8w1pZjupaF2huj2/7utBwg2caonPL9QnFqNhJnw1y8cEijm
U2tA1t1pCHmc/cfMmTL1KVw5knK/j+GUCQdryhHqwEoaWgcU/WsJ66DlhJyiBG8LqQzPrvznCBbb
LaJ3ZRAbBz91jljSVrMpulWLCnotPmY5QRPBNQ==

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="GoWin"
`pragma protect key_keyname="GoWin2016"
`pragma protect key_method="rsa"
`pragma protect key_block
cqAgpvQThUsKP1YQSQ4a4I/shkrWufEhsDBDReUcDIwQgy0J3zK8Xf8BMFoFrewCsS2KNDRzQ+ER
jCDGccgdbKH/8jqChdozG61idZWa0ns7506SogoQlXjlqxzJaYEQMyNxDX7Ycmqi2PkN9cXJyFzV
5txS0QofbL3mzPtdA044rsuP1fkQj0yHft0ysK4zktjTKWnJPMDoc1p9qdrOCvbt1ZBLB18dsflT
y4tm2j7ie4QPZbNefa8AuI4j7gxnCkSCkqJB+CSn4ks4ndlDn/a3c79q59d4UozEclqodJLD4obY
Qe0wLjtJvGaBIVSj8HG9RNO8kRI3GFa3bHt0Iw==

`pragma protect data_keyowner="default-ip-vendor"
`pragma protect data_keyname="default-ip-key"
`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=42000)
`pragma protect data_block
GMWtVErQpQVB3QwSqSu3WLxWBruia83TiqFim1P5yok4XB1LBW9V8dgGNhrpIdx0mL9xCnqViQL9
zzTWSPXPyZIeSD1ylOXk9lVSMYiY5Rh3OqPoNvp3zM3ILnp/zq1QSvEgVe32E0F9UNNyRHxElkDT
D5KCC2YGpVObNXO8uqyNAW/KR2TYC2TUXhdU9vjG+GY5XQIJCygGA7bnKwpw+g6QITAGDVw9P7JA
jPWIW5TM/Cbfx02BGBgwvY4leGcxhsxRUAhhV4/vuHdefaXJu0wXjedwUMeIPYtxA1skiafd0Gg6
78FN8IFSNUOZooK3/yA+V9gQME5wKqC9d4QNxHpsvOO0Z50KnKmYR9yUArxgayzryZz7A6584f2Q
E2lpWLklWiH3pQm/piDUB4yJmnmMJULBAVcvADuK5irbeNvrO4XHgkI20/cer0DcxptBu4d6R4ZM
qG/SfC6fWhVG2lFE7oJ+Qe/3M9amVllSRYbN/dffn4uFVrDmoeaEAf7sf0APiLFZci5vplul7b6f
cSWjn3ZbYO9RtO+J/gnccjfkqGXbVBOESICSXp/Meo2pHJ5Y4NeqdgrUmDVFuTuyiKW7oZBEsHPY
tjcn/ElJpk0B9isrfJn9c7SoMmhbA+d+hJoVHzd06qIvn9DIimXnxgZxQUfRBpAoh5hi00Cbt8gR
hxirQH4gfnlHY+cqpOFAjv94tEInv+IZpNlvJBzlF4RVQvKObf4kD10E/0Xn6UXpOcmQnXec7z2S
JUhwbubAQnduX9FCnJ+8gL0zFswfEJOkUUNpEGsSirEYmFLfXho5g4xItpxVbN6jtiFoQNnIZiaI
4jpoWesezZ6js8hBFT+/m8gc05QIRHwyBJ5A3Y0b+bwA23LlUn3K88zFV8p+re35k6RaO4A4YcX0
VNsEhe7184zF0mhriYAIkAan4S32fSmpMzipuPfWe3ai6CjMIKtCu6oSpv7yFkv91tyAO/CBa+kr
F20ypKWOUZYNZuBNkMn3j9ZoGnEJn1Xzf8XRAKB9Znn+CbwexW/PKLZhPO+rxZm5dpB94gNvbM4E
HtsSq3tRXY4A63l/wmv5K6fJEEmbU0EtM2XF1vJTv1lWBEdjmiJBB83vWCgi5SEXoWShHjGJDxEW
vPQJ3A5A2fUmEmzfLDjnL8REPlJp7b5RuSkCVHScYMy3EFDbvbSQ9/QAtrMVCOJR0HZKK6oZosAB
0D/VcVOidzQwW9f6sBh2zaHNcdPSsYKUox01b4JmF4wyL5KrXK5LvUU+tUTV2Q1mEyNPQsXb/hmK
uSu6L3ZrKFNDCXVMZZ4hoomrOSwLF9X+2LT4VOIBXAjpfwq+ow2Y4CxGjkf+8NVsOutDJtncYKiC
oVcdLAwf2PSDziHsU4uJAVWTjBYv7UnagrBw9TWddMdncF7SjJmmyNpfYrpO4Qphp4TghKY/BiBR
ymPj/KlvuFitv0OhmP2+8ciMpUYVdXUIK1EHESib/ByoJi9FEj4bvGRyoL3UCklLHzOYr+od1utV
OlzQov+UB3P3P89SKriGU9jdDsKZOU3yljr2Jphd05zmNW1F631d+KvnMxvxS85jREoHeBg/ay8T
uvZe57JjTdGvnb9BniPfCcj15PTVCrTygbyWlKFElxeOGfzqEa8KRp3S5440/Ck4EPLO6xLmM1eX
AjSDMcjmVu2Dtg4uhAqKRaBsDRauFy0b26VvBE920lcHgOmvoOsjQRBgXPeGdzWdMTyRxdrPKBq0
6jnoUxTiOcbw7IhIox7PHdVSne+5BOwEDDFIO/IS81sqjPlqwDztFiDmu69T9rm58znnRn/dH+Lt
0xZ7QwqulZGTXbAsEO0pSHrtVA1SC0J133FHm/tDlUm9OJi5gCfm0Hjk3MfvKsF/s7vG2jGJBDiC
Q25eqiYhbAQ1H9cZYVQDUSlrKXGqwmxYzG8t9KHhBLuRMTSBurBdSJxgW+OvDTT1gOeZP8EdQDIp
CDSF/v59hflgcKTqGTDeqhiF7hs39VrCXFFzbOv+07IalT1zj8v8A1wHXHfmj1avRtjRWNkrscNY
jWuo8nwjIM4WQptPQlLT5NbhsGR9Pf1gfq1gHFqYWkgduRs9syqpSSx69AddRLyOZC+1+X2zzS1+
IBGSE/o5zffQoc3rMlc2xChQTBzLgSZl2oAwvlWNixHR+DZCbzjWH0WMmzehK7jE5oPw3S7gU0mR
PFO5tcqVNgApqdRF0xtDscHjMSHyX/vL9NvblTdq3ANqEXOuKZupPabbALt8XQYaMj45MEzFcksD
ZIL1xgAJu4qu3sDDNknZyNB9nufZ58iQqIKDLUvdEv/m275nS4I1Qazue5sEQCJ1ntK+hqb8nevf
Q6gmciNKqB1ahgm9UlbpT+V98l6ZNVgU+YgtbmVQOj+9TA7MnfYtJAOi/cQYTwjLxq65xqw/aHAn
bqRLASQMyrQrcNPBRWoJNbGn9B5SPWBtWi74ucSMFEDU2+A4emOPyqeYXMpD3dYRXgtCuPulRETr
1xJjrjH/vVjsfaGW6t6x0fzGw1We1RiKRLv1K1niuoFutrOJd06ZQEVttT9cvnk1qGC8b1txZbbV
rp4pt4b/TB5FyQx5Hxb0CT9c3FuLN2bVG6KXXPXnN26oFpTv6KeBss46B36/2DKvs+qN2EuFxjb2
FDWin5RddCoBqjCkMFxYMpEntwCMWuUhFv+iYMeeMjOYqUwX9dIZ9ZtAL8iJWIE9bxCGR2hH4z89
qsriuqPZbMJefj0zZMMGXqscQFTuSM7MOXXRfulKrnqtsUrFlEt3doKZZcSPs/ZCeZ4urYmrNjh0
CBvvKaANHPAqH2QEUD4qEcPrEmXMeslqVaiAKBF8o0cICYSn0Bo2HvGCNxLK2C8uJio0fUue6cqL
T205Lgad6kb51pkZwzZJe69hQnilal/mWDg7vDkZs/nITTVGgFlTu+c3DOW6DENlR3C2MOd7dNxh
Y2MgkW+nM4fnunACSYVXz8C08G/dgHM3+cE8NJ8zPsm/SciWusIQB840jinQprGMM5JPobE+9hMu
OEYBtyuqL/QmuAjQnVnzE1QPqd6rsWM4aJ+NyN5lRjDWpKhDc/ra1ngLS5jzOfa7UgNM91/mKMbU
VMu0fFxvNQTeDUo5XaEcCUSDdAWtzs+IstWkw6Ptz3xetvx+QZ/2483ctkPMw44+qD4odxJovLos
eWAo2disgTfKQ0gMS79AV2LbZ/3vrJmvUCdDZsIAYv4dMgqYqWLUEVIUIQYCSXyqSYSx+Dyy4DS1
XMH6j69BWlx566qn9Uk8X1uVeA8QcEDTjmeFJBlxPjAY0B6TDxETb++4/VGEUIGCl2cinKntBOdb
TGPxGJpsLrUASf0F3imACe/aIjTe7HTKJLlrA3H4d9POQ5pBgG2OD+qJV5z81tC91s8OyW9T8lEJ
srsNe9CXyEgJYrxmQLFV2urGh2mnu7wqh9HXpeHRAxKOYFxG1e78+EbdTEfyJuyuX9GavQyIOPR0
cMUuAxotL5CufRMZAv2SgGHAhgGrs8AE75ldnHilI4S0xdXX7Q5DRJDc4bJTvqs2CMIAYYSFiRIm
9OzXTdqMtAKAVUl28CplCqMNJRBvUmUYMN2oDhCo+jYjDbZ40BxxyFjk3pT2HHZYVI2ho4XTXZte
OQfhphy3fm2m+/9yewHQCe8gkN6aoaVxDwVmECT6NQ2L49NKqyKVzFPZ6PG6PjswKUhv/uv2fv4q
uDZqz5RrPGiYrTmF+23DEAJr0gqJP84vgnCT5sdKf3i8HmaCyFxTtkIRuQmjMjgHpBH4yzvhluK8
+tD98GwDqOf/6wtBnBX0OpJq+a1nL37maI2BGwsNkJvy/WTH7tHtYOd4Fo1pwE2hg7my/pNjcT3j
10i76TcAoAebmMtXpBBq2LiiXhng6LM0GKmzsrEy8zv07+DnxC/1PkQVCk6ZyA04Oj6VzRBGxIrL
JUW9MumSrkHqYeIIUqv1aWHYECtp8NQRtWbVQf3B6InSjOJs4nQoZoWceQIkl2hWoULI4JwEVRzd
uZD8yYCgge2WYB9QvVCV+hETpriEtAKbLhH1btyQfuzTCQxYfcyZamoseALcLKdz+9IU2fy8WBoW
CcBm91+8yiAuhBGeMP0liplbkKHGj8oFA9HI7fjo7uyahpuSGurM3yRPi6aO24WzUF2fk+qIJSau
l5iqQ/ONZiOp3FMN6fvPNinzGtl7vmgkGC5q1kv0eJyVaYXqiej43L0BLPFswk41agniIRvuJQKW
fEsKolV4YINBBPgC1sVEeTOfVYdqzU/Lb5a9rXdDItGzKY+CydHMPL5VeRlGEbWu3e/EO9tlf7TE
+SLEX6siLtU/R5i4QNOUrmar3QnA6jgO45fbht2NDuw/LBAgCyReBHxJabGL96w1GlHzwkz5ibJP
bQl4DxWeFD8LGCqWLJbIEOhor339M58rXZpGoi9V4a8ntFq8acW0fYw+3oz8AjW39WQzuaBPBECy
wEWVoIqALm5wn0GXQxAMl6JqQYeGQx4kA6CngiK6WJiQ2n/dVif++R9XUWuTSEDBUhY7D2TnPkAI
18ZEtCt8544rtYBlw2QrdUsMFHTEkf0mmZODGevEd4TnJe6qYhERcyK+ZORLrQKBNliZyBfuM4Lb
CpdNK6DewR2jooIAkygJJMsotq49RBSFGT2R03WczEk4EX8HWE2pHCEisliW6EiDwtYj+Es7j6kw
ORhZ1GXz+BGnKe9Do7zkujGuQMjA+xUHu+sBoGY5YnrJSPztqXDzNDsVSLWJ4Dr8oyiko1L6Loxq
eQKgqLQBQMMN7OvxwS4IsMZRPr60BSyi+mBnFYtB3KWjGMRrXCitSM/PDjdrKk9vqO3z3qmIBK/w
P7043qGEJAq1Q4+8mXPDgOD1eWSx45WUbrESEA8mPcNc1vaHR5eTA5JkFclVCLeg3u/iIM6fvOKq
L5HUY8GCqpWhEqHMw/OO/eC7CTyAYSib5GJZH7ybyBcmePjBRdYIloPYUXhn8uWPk+WfGcguVHWK
OW3f/ceZ+nfJRtb+H5GQr+jo4LEfs+ijpOWg078PYgx9vvu51Fg3sZElWIELKlOm7VFppwQIJKvK
VIozfNAriHz97wbKb//IkHw91TDn3dv407kQqde11lfsOedmdFrsEL1f5ktq0K1BEMTIPB+Wx9Vv
Ve9G31LphSm7TqEZjNoJkM6BlhmPsYB+oe8YSi5xQ2poHv+x4p1GK2lbaAiJvZIgrtWNTIl3gRlA
9Xcan38/oO2eJ2cMxOOIfzW8LsQtWiUh5ZD/PvigvFBJXtIDhEwrSJUvLAVISoz1r4cIAQmGnnxq
vBNRflxn/rWMKDCbkbKrSZwNAy6B5ANo/phhJGjB505YMs8/V8XvP1JCYnIJ7n/2ZPVYK/+NKGTD
PigvDzcT+RqTUcCf14SKN2i+CCeJ53DdmNZF6yX4XQEtBISMV4khsh0ssH9H+I67O/wnyAiSPPD/
gRG7ToMxMCgfHw8TANQxofRixXvZgYg3Grz9iH8jjpP5cm/3ZAF6ErNIrc6XXibNzwmReuPB5lTa
XMAyutRGh5GIJqKRmOcTpMU+uGgtxGAixGBBlCAbsDObFQ8aO1kM8cTIN60v69eDY+NefnPOgEEV
yc1TZeKCQMCC9f7lfqvVx3nK7swgaPxClIbwfPw3XfOM6+l76TRJJLcpT4RJepuHmdb4bRJ3v542
/gjuABa1+epmva4eRbfv92qP519VGC5sM8vxxRLxylNuG0r/SF412gcpHyFzG/AaeWYyeu6yDohG
g/YU8Cm/oCgWOlWwZyhmS37slXY6l8QtP6Inbl2PLAMzR2jINnp+opyjuzI9Z91hThmOxpMmPIHd
4OOgfTVv6tutn5Kkqotr4mxr/KZxBSiR+RH8oNawE4InPIBW3Bgeqo8dpevw1e5mWjoj8SlpSbTr
DXqrfFYWIpjzt0tzn9P7s+qaxiJ40WfvaXnyLnBFY3yVoWgHbQeIabHYcZZ7HghpeEsGxtCvgzpP
K/roMfzp1G811PN8Q7Kpy/43hrRjbkg0TIA63jKECcVdJtgCf25bkVJ40p3xsAD2s4/rgluhOzlM
qZoWl3ZnCAtmBrCCCeMbLt8MqpuO2+hRvN4WvOnuPwWAPRTzQdOxAs7FDpvSmMCUJ+2z6npuzCbJ
HJyDwFviYLcq5YYQW19legwN9vL4DY7eF8AmxVo3dnB4beg4Hdc/1lHXM8DgxeM0t8V7MuweZnfD
3nJ7bJiwM+9fsxnHuQbqM6jjnVxSrEioD6EBVpBKv2vg5RTbVZhE22lUxWH0bO9x3nczejdP946I
13gZtmUhlvSXN1X/agcEZc/mSGZp9HopOBrBkztNkxo24aucQKccOxc8/YblzcXrCFbCqvM1doEl
w6mo+S9GrwBxHuEvX/OmOSRtBe6MWm+lWQdhqReT41T+gpAVpFjl3rQ5Apb7XPf7iv2EDU9TL88u
AO2G+aUba7e/MZyDYE+Ad5zdDD36nW8HQfbuz5EgjEqEr+Q3YnIHFO9x/TUOxH9ooIpieL4BZmIj
l1kdv+1GOtSjlzJHLf6rDvDS+SCgZaCNmIkvwQkEyKv8TjYBWf18ITvb59xTahPI1vgZCMem8gCG
vEor3c9mgI5Sh5bzp41q169Z/HW81IFCw1AqbCnsnvPFhNViD/EGe2S7EUEH/frgxPn3s0vV+D8y
TuPVuDpeFnFxGLU3quuU+CkeMQTF6pxmL9HWvbBrU//nkGFzkT3cizR3SiQRqQQAugBm0qpHmffd
VNlYmfjoP4ptXPHgZ5cuUZWPrgTIAPXpBMajvc7JWzHT89QqoUl1ki1rwDULDQppPq2Y7kR9Hs3h
5YeUTpmDVxCldAiYO5mW8amTzdfZV7tme/NU78kuewuSBfi1S7GzCcYEW9s2ipqMTjrlYJchnEfp
KAcSweOUC4pjmfsgOrg9A6/bXU2NTusPOiBxTWMFy4OsBb+dhxiX76FeDrMEH4LBVb6utkKAEQwU
vvHy8tGJFH1ujJag5NCzhhlDrN3lNXPbSmaGS23KIV/aJMGSrac8ar9JdSesJtaCcO+bRjBJSIEt
ImqdYaHDYBT1FcXJWxmZ59fIzCkenHmedjOrhd1TO/sZU/zs0+A/ERTM8PxphPRf1ogbuqP7L647
A2qgABMaX/wPD1Vtw6iDGwSQxx23JtQ8uah9Ok/yuOjI5Og8H3meS+cx4z9ApEzK1fxmtM5u5KZN
fpmsnJn1vsCph77OEzqYeTE6AzQdXk3RHZGaQdjzuAQmwBP2SoT9AE9+T6sxc837jRQW15EixXaL
6z3bz0zafH7oRLQDrfWsNL6E8vMSk9aUUsIE21v8jXHka6Hh5e9xv1Hm08I7s69n5aU+o6l8p+io
9t4AmuIx1e2BqoGaN2tnkd8O/nsWA823hGPRUbMd2niDEuvRe1K+MlfnrItZ0j/AUIicAXl48Z0J
qJeVVNEBPDIMI3TcgwudTDXgnfBgbnAW29HBdaITwozb1+vaf+0U9DVdfyiw6z86DAdtO2Nzc2zQ
HLkdRM2whZ+NLEhUGScXOTIlpMya6buw3pPFtK/eM4I5tGX1KBYDZbIllbvdfHHU0fNdHE9KhN/q
BU+UuCqPM34SDlAU+7yvcCbecOMpV41eRDdzInlAi/+ZUGZm5RKfgLOcic8jMhZkxxqnQ9tmpxB5
24dxfrsKSwhPNo7EGVUX+0+/8mjQfQQUFnitLpNqC2GqNB9IAw3bY6hc7kva366buTWjFxz2/C1W
S/t0gk/+KgFU+VOeHVBaEasiD9tQk26XeKTAhoDgo2rQ0rIxGd/CDuCj+1j6Mpg8EjZs1HUztM/c
05CzQ6xM/p407CLYBtGYplSlzBBZZ0/wKW3O4yN/TmLitJkUr65ahDDj+OM2t008FyAuwLIEDMKG
BCeKL9XdMJ9tqUIgv5KpAWUH78kUKAOyE9Z35rzZHuYEbz3AUTeU8E0+Kd/5j1qmAtG1Z33D1Aan
KIUdjV5fUGHft51MmKfyYK7tsDQoqOGi55fPJX3eRYEARdEzAGvMDlmzk7icgr1urwjRpL0oUbxg
R0KgUP2RDKKhAKNv4HI/m91nOu5uBWw/e/MsXOMWp0Lv5jgiigv4gPheFng5jE6P0omWYiHU9z1c
rlfxu2g5eTKgcRj431/5chxX4HeT6Ke2tq/5h0Jaw66j0m+/U0+orzrfuzPpjYtYHe4t5KHAhdu+
fR+17OhQWbNszq9WnVasRzDQ5askeTBY/1PxLdu2TBj7nAabTKFVpSk4nkzL7D5FgPBXT08V6JWJ
EpR6u6YaTfj+7DXPe6yXgshmW2UsEYGkAjVKk52u7mfXMP22E0QXue32xH3Up+pros86TAUMWiYa
9TIust242iqxVfB9g9dHqDiDS9oUf/fdRn2dA4unXlXcZJfETx4ptb85GFnj5+uorlIdJTJLmwia
0BBv6P9JjVbLpYeUo21EMCbjjqhTCL5gDSuvsbNmr62xAKfnac7k4etesjjev023SmEgTMUx5wwZ
GBCik7vEZdn0SmUC1d54/YXjoLg7IqITVPpHlgivyxScllZk+WAPI3p+k65C1d2MFBIfSYx57bgr
LZOHc8HRSb0KOgKEw0Wu+sEVLpEFjPCOxtWgSFJdzXd28eRb0n0ZfvQgguIA1tOWetzAoZALoFbk
mME8tRALc6QmI9kLb7n/7qCm90V+o0UFK5Y4oRTeAbLt4GebxBeFwGqIwXM23755JKXPtb6Mf809
2zimvjDC8B9N1yBTNil0+5Y4mlIIbXngO6NcbfOaiGmdd5zvt/6Re8Mu+6gV0+IfGW2nINbo5Uet
WifIy4EAsqbrAwNw3XxjlcrhxpouuBAAMiGEeK9f2VH0HwPcGtdDyOLtg2I/DbgZMqMVXnX15NZ1
NchGv5BhWkAElx9XVi9ceyzzbTgn8AjLoS2x5cGOpPnbJqluEmrvLNz/F9F1M4PMFyd6QfQo3KQR
nwRJxisfz3QRC11K1ilZPswZQ97HAuxTt7BAaPa7BiQLZ7aj1w0gwLSQDIR4YGvTXNaoksTFKpdb
oLT4EiIA/+h3JFBTyAMfn5IJARrpyuTGC75GOmOOxDALJEz3MyWOh2ERGey48AQUsavolnTWRmIE
b/pPTE95PYs9KEVth8eP4WiHe+7kyZxg4B+a9bzEueiD1mPjX/EvQvXY0p7J39XsPtEfBV4RIlXo
Orby8UqLgGAJ9OvQbD+GJWjG1VaaUlVH1qZfGhE3cNZr7mev72nODOQSuI8rrIE3kCHD2JArAzom
fV0WV9s4fmVnQToNUVCo0MzafUhceh9g/aqcN1/4S+Gl0uytL6RpARIZ6SB/4siiXIRDUPWEzASB
kCfj1/Jl5S3TGJ40BMrWN8fI90urf9nmFkrzNn4mnR1AWqyQdIs+fwiBgEgPEHtvDVw0vuIMcH1j
GJM1dIODKxfSRVvwekU9/YqTi/vKeHooSr/idXIo2KsFvdgzm9flo6aag9G7DnAZrxSOpBQ5RNaV
wCFq1eDj1L+rx2OWAP1Fd2hsDvHBLL2YPyGg+kTkXU3vNXIgZi9UW+MpmlNfStdXsLIEFDbZ3HwO
GZFLwYqttQzRpYZREn5jL13HGbquOwyaBKIA3FrewHAovk0TRozij47uP9/oXBeMfVbXFL9c0eJy
wwug78lINoIZ4+KSghooO22Xj9D9JPcTjBccxcSkWyhxodni4Aqlos8euhFNsjE3aCr/hdRCNPN5
QSg3vMTGinfXtyy/wfGOacaJ/mEs9MzmxYTmaaS04tsKbHmaMdC5LJt8vnkNgq7ExE+Zky0ygJVG
fTBwoIJY/ca2E4ymNjbVFIV34n613xl94T60clkUI8m5XKmI1aF1qYQeqzvVi2Xj3hfxq4+vaL0g
zgD2XfrZcJ8MWSsnN0kh1FL2q1uxgVmD0zkdwlGHY+O+N/iEFCGqWxY22pNBxARQ//ML2FSPAci6
TxDYYLQf71oMw/PqStlv511xBks6VKgklJH4D/E5jD/TznmhiEQSscOdqQtefwQoVJXvs4+AawnX
F0I4mvzfXXV24E4f4FxS3NOzQTo6zTcKcTMf1eUV0vtAFI40AgYQuMD/IWsQRlHNVA19hCFxrZ06
q3LjsLOyWJviawbYEoOApPntZjKvRMJBRfb8uI/E59a11E33rR0i5Kp25S8yTvH1CnxLAzFPDdfz
HP1PUPYkTyCT7RJSs5pvDrh0eRLCDBa6Je+N8h0/d7NrW7a+GCeEMhOnyVhusZwZ8xF+kT4y27A+
SOOs/3w/5IHynJNfM4tDiypHHPu8NyJ/Bde/z7pJt+OhBZtUO+AC5Of4E9PcCgt4QDIPANqiclPy
KaDYeoBJLYrOmf+b7s0PvJJDoLDpITjC0xr7xKaqTfMW3XeAAaT7EHuZuipyxn2MdF0b2MtQnVn7
VHFlh6T3TYvBIcut009STv1jimMjVFVZhBg7Db9be8SWmpRo2sioKgYRaQQx1hvcPlEk7TiZUV6D
ZuzCY1PZUrnhBhLCZ617O+sasWlxaH4nPtMY4LEggB5w+aEvYjje3TUBAz9r8lQldxAONAAzibL4
MYnYZaF0e7M3PlWlUl/20OeHzOmvseIT9JLrkVHQ53exRSglxu94RPOk1MrP7fIbsbQ7LHFe6vu7
y5SOSfn3vIptivSeVCencjMar/fSlfSuzf2SvhAUjy+zraHL6ckuayP5LStR5sLaMedU+mcrOHuq
ThRf/hpLRlQnlvKEHuGtG8vD1cZgsT4we9X4EHJ+8yO4yETod8qoyFBeJUxwjllTHWMyTpwUL5rS
UJ7jgknfigst+nI5TzDsq8RFxJY0IwuKEWW7go9iN1rwvyM03kWeM8wSckpvtUWtTMUkNaZ3mzJ1
PTUK30bDAhtWLJlaaS6NPmxCMkVJRLo4GzTOx6xfbBc7k82rgN7uDK2xt4wEe/b3MnjPeQY1BRpP
LM5y46xiQYyWp3XuPMGg259gad/6wxmYo6QCMgi7+I8DqWM2JsvRs7wa3VbwPi5QYAMlGrScu47X
ayx/vRK+uo/CxPirSzFWDFDHrOWiiWny4Nz6R3LJesaa3iUrVEKNcGcAiNeA9McTM61yW73Wc+ID
Dao8hzEMUHFSeLdHC5NnN7o53JAG61SkIX2M4xmtMe/jMWZDCqyN7XimPH+bFq5VxN9ohBBE/KhE
u00gaG6+TYzKtcG9edZdMlokfhI5maqzP7Y++GObtYFHfKIp3AaYCLw0BHMTaSwCKQbbrtTnIFN8
6A5enl9ECBBJk9xFwxHfMUeZDlfmi8Rdr06ynBGvJ+zuEsUjjruLdBN65SPqAWeNJOQ9aue3fBsM
xvNy7ll+/+bbF6KOF/mYDKOblORKi4xT5T4WNy4W+PX+OlnndYqX4sRPfZi9b5fWU/ODVWZuPUZB
hKZ7RWVXd0a3smvqRyRyHsoY5H63PQuk24g7y38XG/M2ogHC6hnK/eWK45/UNI7UFnccCrntcAHM
dHA2qI0kEkQ3SCwAunhwlWQ7rFZIDbJzE/KtJgl3K6I8quHlaXPHjPorrOp+YBnEaZRvW86MKE+4
NSOLLl/L+JmrMLI1GdijPO0PxGkG7mlo2dq7+Wz/XirsfjgyR5qVvSlu0EbU5172Svk5lRjkfMiQ
bb2gG2pVjwDIMXyVkNOQMMTJUcebcqYuqGKY8papzDe10iEx3bR4FbRlJNfSMPuQxNFy9+35tsQz
UkDeIWtcoU+Ls4+d9Ad4YVavP2S8OArrptbkrxGKVLhhat9cDPIQX4+8tIBtsphOlA2EEDa/glxv
890StQGiQV4a83bdVq5klwp51WuQH+56jbKQlmLujMvQrEB92LaDjQfBG2U7IGppQd0ROrVLbrel
MD8wfj9hpisJqvTjoi4rtVE7/olXOreYJG20TVyYA1uOyRf5fqDgE3erId0EaEfy/z1EWrCviH0T
zd07EKoZx0Xy53mhxJZN6f3Egp8nHgA5KLu91woa6sQw1ZRURXPVV/4T9IFktnwO0ZbWRZevK25q
Oqd06YJ67aXV8PEsHi5nUhmvHX4mSt2gt7fIZQ0BRbFKbSMWaDF9185zoYrSkp73rMQzMNN6HgQ2
HmEV9rC4oFJuOQJo+Np0aghxPBUKVPqoODgX3rDFm03n9ibYskF01CGG2xS5vIYcVqPNftxZEDD5
gPQoNgE1wMQNGqOg7p91ai9Tp5vX4WgrH+7MbJi0t7s/u9ruDQ+EdVH5U5VqQDzEsAJqrK354AbC
yPJheQraEXSH0P6kdwQxFpC+zRXoKo92Xi2DfqnC95/OeceQbaakEYccu00h9lemFN7Ap93Pt786
8XXeXF9cM5RV8rFKsFzOAn9yI34mwn/vXXHunMI9gFKpuhPgIqoIH8WsXjZ4lEfHLXr1fY3CKMGN
9UrXVBxkKQdlTg37SV3go6r59aBaaVkMg3nGiST5zmueZjwAci2QcOIrLiPQGY3DAvpydu5E7FFQ
jeLwDvGsig0Kw4FqnlB4b7aM6dpspiMQH6z2p6xbCNdn3eOh4ry8zwwhwN54qZEZ+FjVQsfgNIFU
mVsXeTVHeIWETVSTIZHWRLaFJj2D2YgVZGYE+w/LnNA3ctu1YO36xcAHNDs9oT02aZgrqzRO1Wqn
DiJYBFWVFcLh3/Am31vqa5eBP4cKT/cHPU7y4tDkAuLyhwzXVSnD3fmgArEzErvY6d0xh9oY4Gpm
AxhzTjh/MNtAqdIwXKGEaAlHp7JtUsd4rEKxyflCZJhPcQ/ZN8AC+jUyoeuzw80lOtlED0dTjeab
NsH96CLNDkf5QbMqFohSZHw6SQ+FveMLt5YwFncSbsYfhFa4mJ7x351yAPBLuS2nEIW0mLlm7WSk
XULzv8eQp1NhxNKvqz8/jc8JCcYPl9qDoEtY3csLL6GW8BXh51nUa69qThtawAWbcrzTPbDf4wfo
P2iUNHUbv2eUlZr7jRAKfu6d0tRWaUW3NoAiV+mz3D3yRP5Q/Rv04Lk3lgA1dV8riXcgpJLHcRt/
nx7JIwShaxF1J7pHF9EM+DSpL8XjAa9fHpHCYPvwPXwm9fKWTYjqDnSz5//KTQK27JH9mw8ELa5U
BdJbFnrEQyFtqvGSZViqjoClO+YA8ku72TFWSbnkP3FLnIUIfAwsHwLzrC7h3zliyWRN98u7+qEa
MwLthXXDGq5BqD/kwD4DlYytM1yVdQTWMMj/zvJcmeniZyM3EmkYYxMa+OXkUSdRTyTk+2k6zVtP
kyaIz50c/Xje/g3Xj9eqaMnQ3R3zacRWxEcMoMqyXZ2sKLZdFtSVaVTz/4BHJM9cfY/8K1sMk2Oa
jgT4wNC/cIqi7GAoKGDeKB2OkAYGkdSNKImid5sddMre0kjj2+h6tCRlbIC9D12pmNeP0bwg5ojS
BzitQFXLtXv7nRVwWUZ1kA9VMI9oWD2jYJfpdCrVUXlU94BJfmJmFHoR0o+49SkPGQDX9VbCaFE2
uEZENPApWGcbXmEoITjk8NtIl5cWm3VYU+P7BjNK99wvYU77rObw4hVpcqumhLVJBFX3dOBu7vXD
IpasxDQUvfddo7J+KeQeNUnF1dxBtOjRPNHTJzpLP7/5SaAYy2emwFrS04vlM9YuZTMjx8TConqv
pSJQg1HWzL9kZjwEeJXO5Z1MOeLYKlQCaRtiUu4FG1DS23QoHMEG47hk8AFJ+bNOlm9MbWCE0iFr
ECotw96uhSUW+5On51j5IttPeIcCR7+bEUR+C+WIv3OU/7LVxva5GRz+h52MrmZ+uKAG+N0RgUQx
kQxd++7DUqhdBXhZo8nh/m6j/bl3Jus61ky21JYLrNrTdt4VnDaYfruQaRo9iEAB5kmJvsh62EMI
AOFVTonCm1n4gwtqsn4eEPlj6di45AOV635MktEsJ2TfYvyQgn71imcBPveTEANyEHP4I20O/5qD
L+db8R/aU1wvVnhMu2p326wGnqXGO2DYRJSsnzm4Jj3KLYA3mQ0Nd+kkBE+GG5LRsEh+2cVsYtIO
YvqSBa6QWEMoPDJKHy/UYJBwaLj7eu8bkdyGmvIrok8pr2j20FPw4uFfDl4NF9+e4ArHsBML+iBR
z10Sy4cCZkxicv5BjtXsDntaeOqhIxju3dKZiZeM8n66CezqD/jkmryybA54MSO1ooMC0t1bCBxU
HMJOeURX1M2FVuw4+Jrw/HKm+KNGT7t7uO/4v7+HOtLeBU5TJpvS/ALFfTMu8/Ub8G0Y6AN/wMOl
s7ye/Gl5LQWCC/eVcAlpw2RWRcu5+xUMYTncMRXk05flzCG7+qzxh8vvMyGoYg3YvOPIx8r0hATN
SuMfdcKUxsEwgecQVcVYIRP10Defa+5V6MaxBQjbUGj7GqiLbxjdYcP3jyrtfFcowHx4XLitpn0+
RONoJbPqulzWZB7Bfm7l1pIuza0qqk4KTymtrUk2V8nQjccu9aMvajpqdCAfl6SGZhTCnSQxx53q
9zWPiF0CrrEd+UZdEpCXaS7uVsxO0zoeyMabJ5TT6iquYalSxACRtvLDpYusNi+Hqj16CPkaNzeS
FZ0f6qneAx6vZl51wvk+N4mOklVjyUEGfnci9/eDqP9X8dUTeysiWRoJw8ZamC3ThI0Cu2Sn7gju
SGg9dZb/htH/zblS2e24YNJp+9EptE1B+Nj5gaeOBa2KLbjV2fV+VJ5VyQ3WGGfiiT2Wkf7+LMrd
eeNhQME8jazRg+5kAcZGsTXD38UQ14qNYrhWNc4gWdcfDn221L7cMNPbngkMGGN4br/l4uq/qetX
Z6Ly9DrfPF05aPA+vOdc2fDzqRn13pGU2dgKSWDa8MVRqf2Ry6BaAFcOj3nAjG2shmdLjgxg0xoo
1JuaiRZsaGeQo5k/QKg/Is1xfvKKdtZJkY2orLvqSNlR8PWTsuJgQHS2kw3v9jeh+IDw3GcdWU5O
W5SjuxOcSQFlk4+DC36wOMvyBhFPEnv0yiUHLl54vVH9g8cy93K0OzGWt+w2sN86iNxgmU/WWSBH
BBuNxPsDcm+fxTibSo3oLMtLbdbHcbakW4L/UDc4xUI17/qe0DKUS0rG4OgD6U50wuYzA9N+SqSB
UNfotTY8rYctmAmoj0omrefYbDDDk45ubOBl8JuD2agMfFHne5IrfjWh/VYG6QXCFPf3QkX5DbxT
xVGYRC5Ygm6yae5p8hyMx9W95eQKymm/vC9lSKvs+edWYHNnlal8v/HJzdzKi5XX80R2m3mqmuGq
WEsPUGWw/HAHuauyzCH4KSscHge3oY5eRVsb4DdpfIY0D68rEzIfgJPtKae5ZPux6ASDLCwTGSqz
j2rMIDF3VFzFucqGZPqMfb9jH+BuCIaWUkL7ZyVxo9wQpchPwaKW3uzJJxoh8NnmsojSDQZWoNa/
wZzx/hVh7SZkhJ1l5sMYJyPgzI/1fC4/Rq5+F4vQkH8eQ4ASocxmWUiZtGq0SfA+w7bJeqC15Txc
xi7hzaRG7Iin6IClwdxRhwbq/Le9VJ43OOArNG9B6Q5jCSvp1sZZlnx2rA/SFro3Xlpra6xU09qc
pcgOSrcBO3Un/ix1b0o3W134Clz9gNceSYNuiu0rLR7MTwJOGMox8ZLg/iQs7RhYdDwzSR8euPiM
zbm+rdXosqm9rZaEUHaUy9sr2Vat6npvafHPSmALSfmqOwyvNUtMigwu35ZdyE12gIFfBxxX5jth
H6YRs4SgA5oRERBXzpTW4RMswSSMO7mrQoJA1dJCPEGcs/fxUJpH2VroQEG7qkdanRuOQEpb++aW
8a1gHp72Bi5fxR5y6RdoJVTxDcq98XhR3Ei/ZtmTzd6M6q75NEzuQ/lhziTckCB8qLH/pWVfvBPE
/LHMWSpbbDKXnlCJGTHkHK/y518Oa6r/WLOgTZ61aslRxiKPyN5M6TnkOVMpIBP8LWt0PDjwwge8
V9p/K+MX92Yhuh2KXC7/+CCT4kq6Kpk2pEiQoIKnZHJpNBA6d2qMG/i8pNugfdaFtzVuR7X8jRTT
NrWegRwTYLyBUU0rIXeds1wQb1udmki7zBjC+aE6IqMmzqPaPA/P/f8VYaEWEP3HxrdoVtlkoxTY
rZp93pPvDm8wWmQHphKk1coixyC3OhPSjdWAQ6N5RFhimw+Mc5pFD+oMkcI3Y3+v64EAsSyOMhBP
pNlNA6FiG6kA+SeXzxaY8OxQikZLMpImNAal2K/V+YQrpoeBRgnjVhEa+tLIUvrELUJbo3ms9oLr
CopqtzTc78aT+E8yjV7tBL3WhlonRcaFpiKfcjHGy0nfMlDZB5ZH5ngmLmS7+I4v8uutyeu4xpck
HmNvIkgFC1xtlR0/dlTNPN+H4srAcoG16RlbampOR4B3qqYxmVSZndZrtw78VjIvk1SOSaxovlzf
3fzzw83qzkiCY7LDrhkGO/fdWCdcSm3TtPVUWc5hF0j1UxIfOOO/pRsO/4Mw6bTR9lCdBVo6wRAy
K7MsXQ12MFJoOUWiq0aJ/Z4CXEzfxwgjG9Sopq+px/icEqozpRfEI3BANYQD1LBxuA4AeDBuvRqq
1cfy1/UtvZDfnhs9kimjM2RYbS35PZ824Q7k3ZbXDQpLp39yhE7Q5tPjhPoTJUCO9MsqRv8JEXkR
lh2Fu5uR5ptSUgNsp1aMC9Y1m1m4kaBhtCERp9q7xFl8piconpcoxCP/p7yNpZhRbmXaf9DN4a03
Uv4e9iMwNbZ5MHo9X1OvQq6lV6FjlTl752OjH3jf8fEZSpP4DpB6byI8S3rZsZnLAowUXZ7pdzpd
SPqpcUDrk7fGqYct3kiQgMT5Ai+iTERVwg+fj/NG6h3xTWBrxJ6u+aYMEVPydXDNZ2iOvGY/TYSc
CTlKW9LRN10Fgx2QbABMyEv6dGlDmGCiMEZM4nO6ILejED2w1co9lVDezC5iICu7hLEU+IhJR+aQ
RPioIChVq23Y2ywS/Lhx127emjA9ST8Ti4vVvHnwGNpVmJtQSuUWcf1X8h03hWJSTB2786NMSpTo
c9aBjZBa1nOqzUGiYH3He0bN1adk1mmpi8uvR/qezV5boLMMo2Dc1aNTP/NLQNvoBNjYYV/LvFdL
BHAmOEehxxIGklkviWrLUEqoGAbxiLf+g9ajTnZwYF6V00T2sAuwVSUKWNVzV1rLBv5h8AyXZg5f
GXvL5bXy+WiBQnvPPoCRwnFRKas4QzwaZ+lr0JrE+Zp8qrXDlKXRgpJtpQwHmO1LwKdshwUv+GCc
o0VqHqZDtuGRdWEnmpoGCyTaHNrdYzBYT8PbEKVZIl6uy91YaL6ilAdDD17YC+YSzTgD2ThiAKat
dOJPE5b9UZ9jFJ+/epkYXJhwaYtubWAcGs9+7HwibFEjfFPBGikLMHeRU5c7vMYL2joWMSVaBcju
2s8ECQyYjHC+KRdJTA344N+Nz+l5s82cM5mZXu/a3ewXiXSliiW1AUHNzkeEYFVENF5fubrWdiu4
StJswm+Ji/1Br5KeKq0jXoHXg6tEtZfcPAg7PZhq1T/izHKd0VfpbiG3FbHXcUYXts0gWMAefxhV
1eHtW3jrnoI7VGwU0arzndMheOBhLnezUjs2p5WiaagyUP6b4v4zNxXdufOB0nQ5TzA/CaCr2LZV
R0YnPylgWQVRJse/zUd6LTmw9c28uvia1MkEp+EDZihLuqoCE3uvqO36iQ8coFq8tFtbuOxFRc1U
yqNK81cfh0QZEQr0DlI0PF9UfylKCj9megD7Bw9YxueGyg4PgNsyD12WZEMm57JTu8dwJcPOD3HY
7GBwpP0Txi5S95Z8ghbAWi05V2GYk1ltQdjJQ9wV6v7zaEBYIEfWqhNi7RYdELepXxnKRyA/rxEg
2U4wJ2TpT3TDOTeusuHpTxCFxhv49KY447oHqYLDN7RB4E/HSQ6nkBg7XirEQGHwm0YxS5cM0kLa
IUlgrjdNd+MF02bv4uOjnPWcjv9QZWQ8FVYsAN5R4ibv0H7juC5aC9ecRFHwAr7XJbXjUs+hHR3j
9g+vzKVIf0xkoiYztaKEbcFG4m/O5w6SnTKIBl8IvfI0el0ezmbW3AhRg8YHN8W6DPsPJwDO+dP9
z7TX8+o/w+QEqyn2VzGGCcNY3bCjISRvUMTfz8fend3i2El0c6f+Ax7uXINVmOluaBsmqzq4q57u
ptwO/osMMWNhk0UE3wO9FcapnbOf5wE8Mnz1zF2eec5iCFVcZQjRh06t80rstfS5vgqCEFiacHDP
V9/rLAK00cQWH9rrQXCJMQVkTOoXM/hiqzBPW20iBdtPyHPAnRRyVibarEVNK/hpfkmS8+tuIWy8
Hz8Gl0BgBE5L4yzfEZ2oH4tPBQtlbZcLETOYM0ViUcO7I/kd7zUT0fTaeRxlrE1OSyJbF91HchZN
C87mkmYJiAQp3jCYXWjWh1FMoZ9I7omWvcrCx8L9fHI7hSJxXtJ1qbxvg/CqhwY9Duw/7EBfY55d
3mrG1Ilu7MkuE8tC/s393LLnYPPwxsY0efBj6sahnqPvDAsFs07nINth8nmyykIKXmPDqQz399NH
IwTYTdrQmkyg/xAAWprcMnE9RtMW08zMwxpY1wG+M0A9fLfI3Oj08WCEN/adOL/NcBmUQdBnngB8
WIIUgJO3lAOMOCHnoMTI8KAcN/rDyEwkcJ4ogAPHmGhEdvtr2McITJjr1LbDgYQtZhs8h/rgbASY
d2542NvvtTCs9esiDFt7UUrsL+2ngjdDGlBvM+zb8HlPeQY9gGTl3zxYOhEUs6LXCFm96hzQ/5TH
m9fHkwICw5OQmJHG59a8oS++kfiXjfyOAhrIVZbMtMtT52h1GcsKQJ0+ZAKOrNj1C9KmIBt+ICfi
itU/i1/B1gE4iysAsw0ttIuyzpD7iBIwFWshml3FxMX+YyGwkiOTO11EFj16Kze/K9QoQ/tuLO6Q
ouy6lN6PZ7yX3lZ4TdK94ERQNFf6ImwsadT6c4meWLgubJQ+GJmJK20MTjdRQVGMRQSHxXG6BY3s
LMUvNI+L9vFVdL7c3MjqAlcbL7hinN608ngAEEjasbrQv2FfHV2cGlL509i08JtGuZ8qmXbjtbxB
1naE7XjWF5F5NnkUCIDseWl/ieXrbQB6+gpedr+awoL93+/7agqm9XNpzp69eBVc02hj4Z6I+E7T
kK6LylYoYgBklGebiT9TudDcHgxED3Qmuu3sxuz/1n2pYaQcuTMkkZWNVjGYIfYt/cWOK12oJ1eg
UNSkqidiTzc3wuD7ho3LDpal4KFLFj+9+CuBf2DxW59wEqc1dQ/w34ifTYdjTtJwEoXArzGq0bqX
TYjTLixPZc0ldD1JsuZkPxplH80XmpGGKtO/zxO/CxUXdqhajNOLdyaT8SvAFFs1rl33u0nqBSLU
Mo2po18VZ7ZL9dlpHgPehy5+QMGTEUUMrYO/G1nCmcXL2tU4UpBXtaiAwKLBTU22p/pohSYkYf2s
/4MbFd6VZewfJ8Sd5pecscw8Kznl+25OQhRzJuZ3dGwbHiFVAV3Mdr5Xy71MjWYnnjMAas2eD5xW
v/KR1ypelkStDb93mk4FLq/9M8X/lkdAifmrqIa8vcZKS7utrPV/A85kr7jBLKMEUu070r4lmrmr
q3NRwxnLxZa1FFmd8oNHtQvjt+aJzWL8p+4seapeqM7hXhnEI3rWxGuANU6Ij44TQR7aZAAS7Opu
3ueKcxiAXkEr1AZi+STq5Hta9dqFiinnY5BOYQzbJDQLGO/7JhTu8FuYCHhsG3ZtICrlL2Z/hS+m
r/iIQmjzNeD+XE4sRccfKbOB7zK0W/4lpg026GPwXSqtr3UgLELFh0I3nQkmrAe7Hz/Zjj5Jztmw
SuAcxHzVjLFDzQ9OHABUfBZjGwKymD5WwGe3v9RAo5NZx+kl4cwFILGBMySfu5USa6QF/qYLTr1L
Em+5WUQqvYLgUHEeanq3/ytr8a4HNHO92gbCpAUOf/sDSInkuWc/NOhnjGf4Qx5cKMvIm2fJnZOy
31grs79YMv285I+VqquRGUOObc5B5+EXMSjOCLReHrhHvTUCoJlOglC3687Lzda0jYDLZilzCHrs
XGFSOt+DjAQw1Zironp15Fga5R19Bn+vNo2/vHhBk+Pjzt+jHAAcZ/j4LVmt3EoapMKzDz4X5f7F
hHwlebRTqyhq5gAbUazagohm/2l9+WpWveAypzavbIasvprv6UvDKOvryNShnahEXajPbYWLG0Dc
qagIlWLHO5O/E2sfQF6E1IVFoChSCewCsTmoaOj9ompPzbM6i5jctnOzzhGGbI69UjELsJ198viK
ySpER9skdseF2qc05p/fUu63g96ZTttXdkWeiSuEAGDXUOsovOjnVM/WfK/IOL0jTiU5MThlM/CQ
q5QBlvBgNPRGI3TIMTzQ0HkVGNsq31qPIzHTY78aPwnJ8nMMbU+eV8YQ51AUweNwMiByTHyJNamC
spzZOaYfV+zHZLNGcGyNVgccR+eumyyOf2jBrBxjzDlKNJv007LwuxIF0ozMlR/n4LPm0EE8ucK8
+b2Rchkvzb7TmkbBDRu7M/w21qTbt0TMtaTbv9no3zEvDpYzpl+p9QDFlO1laebwFZ6O1DjUgNgY
ejM6+AUUs8Y0DegjWGNe463nkQIYkdbVLVmYfn8lcPX6SPEmZ8rP3vAvB+NoRVoaGYo8AKXenxqf
X5lyVIX7F6lIDgDnxBTAgpteOW6C+W3DlU939QcLVKpns3lA2FHqkNlkBPg9FNLdFyi2IRf4VH9X
1FzVckkOf3SQm7u8yph1OW5cSa382tNubR879uuW+QIcDqEne43YnjbasnVOTuQVraqvqYlI0wAW
MBc1LCnOEE+BsDRR77HMsIf6OOMKPzsaeQWIW3Z0dqB8FJCvK15z0rULYFvFvg8dwXBQviSFgk9T
+b2FScqPA8lFB27OA6sczmwW3U714Lqh1wnN0tM3umhLvhgs7KfH37heWPu0CPK2UmBcHfnulDky
N3wEYtJ9UEGVxwkAV4jZv5PwYN8EEqwm91D3F6gYb7WvB3ytpmTTts1cuP4ujJcghOOn1fhrYgiZ
7uVhQ4QOMVp8LscnnyiRB5FS4LihTAtHNg6hEmjNbQ2dgx2waGeqIwGGfcKgAckzd8S5tl1dyswq
uRyEiFjgC2kSAg6jWdSYKDF6J0S9Q6Zq/V6Xp23U66OLullmqH/Ui9KIxxGNEgHtWY54JrUkobbH
FQiBn3VcMFsHfBXF5HSsNK2ChO2WcR3ov5VyN+gpvvnFyUFi/qAFgPhlZPFcoKuv47djZGTa4kaN
frZFm0vXhbA6LxfWHS37egfm6WLmulyd7H6ryinPFs7eRLFR7gVQN8PITxnYvfE48SZShJ7aabAP
+Dp1YP2CGyW3NKmdHsfrzTybS0MyePHA5khFdYdRoEdm5GvWJzwk/YwWBhVzycdyq0YZZJ2PWczv
moHubuXIaQud3VTN7U9u1rS2Sh92H52Au6AnSJwhRaJ0I1ne/DQK8BTVWIJ7jXZ6Kfe/IZnnO9ds
KJ1tM6zCJRrA0mY8mKEXEHZ0reXTj1LntTtyMgwSIehtSPhfzeC3VMn1VxzKIS36PvQQodhWErpu
KEA1oJcB/0L4ojjHO5P079X8N93o9HAcxl1YpBZ4oyXyEGgnaufFRIkFTkqaNLhrzduXgFBEFd9P
MALW8GBu6ljBRa2NNJsh1eml9rIyqcQditLZfWPEqQEOAHrIhjmNhessQlYpLItLoJsROqiKu1qK
YrH7GeelG6905qiD9lVicbksWAuI6V+EHJeLwajQX2vjytQltgr2RMuxx8QMPkeqQCx8bNSHMdx3
Y8/UZ2Lxl7L78yPXxO7ToU8oIW4XTbevqQueqO7C8TuM3iJODjq/jxJ51pS2PnD25yQuEMBgA+8i
OO5HY/HNB3cZMyj/hsSr/HBw2O1Tyjq4yRLnXafgox9ZuqvqMohofmt9fEv+csbypvEOrZDZb4vX
861mQa3LURymIoi+udln+Qvxxpf7WagO/WSO5V24App3LhRLYUvGo6DcjS4wOZClW90dqHbfTy0D
gRFIYMdz3vNSN+ZTDKtat6wKxx7gmaGGKCFW6QdM9D8xZe8jRRes5WmCgYiH1etCw4Qah4gMK6Lh
Og1/Cw35g3u7Xg21rhKe8jvJ/f/+kf3BMeO4YwnPY2BkpW76V3JS+iAdtssbBSqSi+yKz9kmqKZX
IMC/HQuXp61vEI1naqQEa5dZwqbf2EsTrZnnz5ZxtWC6Y7VzurTG6uh3tpWAj29xo2PdqiM8pIBf
Eg/G+IOBgsY9d26f75165HMMFnsxBAcRjQcZRRAld1pTrxE/jvT5AS731v7g/XLcVohIfkFcpeHV
3cAP7ZQixFtPa+CO0yOrusIFA3tmZBplhKQQIV5cZQfQH5+fahmWN/6kX9NMsqoOMPpd9ix+ys+r
4uISGDyWlcCkEYfuXoWHN+bmR3RnScBU2kVOI0yadxdglTWiTuwndqjAV7uPgYCOCSwVLIDus9ao
TxWT3ziG/7FllG9VQZdEojDQHKmbT/atECuifwoTTyQBZmHAlWjIis+jVCzroBOaNC/1nBhyJo8L
4fRam5WOhVsi/xSc7pm1gS/5PSJXM/Soc7EZxYO4tziOSVxxva/u1kIrVFSvByU5qgbYpeqS5n3g
RqZ1pFolTJo9OmsppUu6PuxXnhpWzrymcrd8FB0gdwc6p6ZoggYSrvratzJuUDHJ+ROVWvoCtqTx
pizwMxVdcADdcDQfJlGMP8wf8FvVZbxiLsKXl15RJrL3cSXFNVXiqDacAYkWQk21qMRCWRYwi2q+
PcNAhBcm/NdeqJhemOmAfOYS3Vi6hCQr+G/ZJrI2fgN5qUtTX7kR9z6o0abi88dKRNJdGwuSg7Ub
+A8RuDvNSkM8w8se8xQMrNTKD+czep5fLzwyTPTDnj/W59s/7HdLec3rwog6GW9px1PogwkAS5/Y
OYCxwUcUbeuDn8hHSinxUy/b8kRU/ddjSWVubNkprf6v2HBFWtEGC/02pZ+NDfhchVjrzvS+JSpe
zb6c6oyYa29sz/H3fWzRJL+PzxLjgf4TLEmHWYfRCmAYLIu17DRiz8GEi8loWPR4PMF9m+PjJ8nx
A57OiSZUI+anSA0PMXtZRNWqfTqTAFs7PrgTxnmRDr1a9FC2Omw85D1QYNw47o5YMJ/kaziRvKgK
QwFXXP+Hl31n47Zwn//soKJH0j68Qu9SLpdI3GbmrIYlxOVGQQ4UOufq/oUsm0eab1jtOh0Xc7kZ
RVaZAxiV69SvSCl+uNXSu9jRfsJ2jorVGU5voXZYyElHS7Wh5+1gtP4fzTMeuefgtYihyMbs9/7W
6or/k2Zv31CiISLwjxNg9wZUVnS75oEjGv7OHSGHvHLEhFNWYhHudaSgXgSv6X2XEHAsBKQ9uVRU
9/F0tzl2stLGUtehNshCTynMP5o+Y1a8kVnzf9T/wXWNg6pzgIlqDXZpRRX8FTxLe6tBj9UFiixo
KtzwUlOVzlt6CjUFsTldP+cGBfunL5+l4td8dLdHxOoAglQ+tGuX7zxBjVlMvPbkFBMnhQoz6CNb
jJceCsdASo05mnutZruokbldr0gjfM+BvKW0CDTzUoY9ssrhEKK+dmpFEH3BT2LF4HzQrfnaHbnU
oVnyMSdMGbn/rQYK2ZMXMvz5duhuxbk5ZZdVPfADA8WMYDhZZbLhKf1SAetyNcR/mXg+O9CDlPvH
a3U8sNDPzq5rjEZtxDY9aPImYgIXVfNFXLfAJtkvYx0Ar77dEYgHBG/oyZhbKdZfAd1TAUFLa2cK
w1oKy4RpSyjB+fpdjO0oDrrtZC4CyQ3FbWGHABI6m5lVyd6NRJp/d4aP1a7tCNq7cEX3naa3HEO5
MmXhlcT/WPyni1oSNH+6t6cQM8FK5gbXtQUkLAeBx21io3odiY5II3NkVKaXGXSiulTsx31hEJwo
C4UfsLEZhF41b8SWc3pHmvGLJ8wcNP00YqopNZU+9y3P+A/mr8ru8n0sPXWckiPjYFCxSpI6hrC9
MlxqApr3HdmgBziwc5sPFdgL5a9fKLmnruKfpeUXn2nv0kXRglYgc4UuLcw3mlXIW5GWLbFY8OaA
DveT3l2APTMp9Q16jXl9OCCqLqB6CRIMbxV2WLPYM1kdMJp//HUmd+e7tx59gqso93cOKpxGRX8T
/ikqOvY7FOVJsXztNrhoGPKKp6MnIO1w5tskJZvzT93m3pu96cQQN0qaRqpCRhNAnMSm25bI298e
sbOEUuDFPk2ooVzwAJMIiRBWaiBqP0fkGjXAZ4+LcocA/3mQiPq24+k5ZStOr3G8+z3PDPtOPFBg
ru2TLtw9VyvCJA3Ac+eXvDRSvCXheb0O3zIMgZhW36HsRez3NsK2stnXu4+px2mOmqjdRWPhEsyr
Pm5vYvDuKoSKavjU2TxuvpGUyhhoMioACgFGvKDv7VBQFRSv1rqygQkA9N1XDqrcU+w3dLNLXbv5
dKvy3Dsqa6bz0uQQs60Wj65Du9iiLE2Bu8Qwn8eJriUTgM5fiChI3VYo91yGaUwXFbWW3s6Hf06C
CBDaTHv5zaGh0/YSSGs20yCHd1QeO0VnxNPFadZXtjRWNiRk6xWmZ7m/pSH2iCOFLWrcNh2KpTkK
T4cVWLf7A3JMwVG7dZ8js8UyhhUjO7YILxKSjqNL0ydLy2Q62lsIMT5f5ru+TBXlli5BweF/QHxG
wLRIs3VWJTefZe/wp0crb/l2biT5lh1xPRbp9oUHseNYCzcE/sSHFqOnP5Y4Rl0vfYutn1952MoE
jEdK3PA6IMI4xis6c9Ck4G59FU4RrcQVWHdpqmCtGsVKq0C3zMQceA+s+/y93ErQ9tujv6JuVj5N
McyzC8hgAdchkiM18mlaQ8VC2SlfvYMjtxHqZsTrEjAW/0MjcJTQaw6DmFgwvCHly0UvwGdfBHMA
xqz23LeohSzbRYquhXg9Sm2s+5WXL8SMpz7/X8RrUu9MuFUJWjy8gli8ozI0ZXV7El4gY1Ek6BrE
ejy3pf4J7yLvK4N8zsrDk2c9naHEuB9r2Hv0loAe7cpcx3rlT+kYinH8oWR5WU8mqFWdN/0h0z/Q
3kqarsFpV8JRoGkvD6co4C0qwyN6SHSP3GHgrgOWFeLOo4pqSxsJh412GPaJGH7xsreSzei4QgcH
EFGjBu4kSTAOiVLEagUV2YYBgb72XbZ8EuySqD1KxAeIDt3bW7ZalXxNWU8uodQPmEyMx4fl4UcJ
KKzme6g7jko9YURgDNpwexGIypey7SO9MotonZERSAs73hs73Mf91ZNFPNjBTCkL3P7niV2uA/hi
I4FwtyvEdmr/+sAhw1mErvPBqVpKoAp8bguYmH2tXQaJH7BI0gljM75VHX551QoKBFyO9S/P5SSe
D9dRzQ0I7r2ULR1YI7/KwToDIWzagUkGM/QDRqpK4uw7Cb1vSxidpAtL+fxEU91GzBlddHOJ4GWd
NQlJ422WVhP9ALv3ootYtlw1DsUjafDx/jogJT0+fv0FexLLlGWJxvJyi9oar3CQfRxqeNQi6VSZ
QVLnl5MjdkigrAQmoYfettV1MdJY5z0Yyt55AaBn4xoJfd9r2RdgXFcq/gG+nf5dCudqdCmW5ca4
wV5vdYhJx1lEmFdBU/jEqzF1b0gNJfW4yve1aKq3RfFg5EbinUVR9DCmcSMHWqOjDeJqEXwDY0Xg
folTcMhLRCit8o8dk9AjBlu0ZKfGl88aMrYctWfWzVfATNDSQe5bzVc9Xz+tvRMRi/MAnWuaqHbx
8gEx9S8sLWMPQ8PvQduP27oNCDC5mxR85rwao2kTQ3FYb6A8lyogRr6GvTA0SQjz0xak3XaLUOXh
5VyQuVv0wAy+kYtkyDkMbGJaOAdESWgaDt0rOnp8fw+zwe42J1YrvUsNQQT1tTsYd9LHO7qCo9ow
AWQm8ZNFYKWAOrm5kw35IkjhTYr7r9jneUYqj3RFE+gyv9CqoS9fzb1wTMIeoq3IDPj0nX1buTly
zgOvNCHaNnDZV2wPe9y1+OuZspD5Ua655Q8Aat8eZo/V6fHrGOb9yTV6sKay89Q25UlRLrpPse+K
wYmPdPn6knefUjXnxy2FQSKq9uqOxtubT/bpWvMjxtO4AO83hVQTEiCgyqoWQJKUSa/S9XFYHpv1
K/UIFz8u6Ru0POj4o/sJRs6fbjQ6ci8McLMfXyL8QFfHnXoYIUYs7Ftjmm6TJMuB4fFmh+cUZLJ5
xAYDwoAVPk9ZI/K1k5zJDuEf53M+V6MJqdelX7BHG0HrYkMiAtQZ1aDjLyHPjOa4cjn+ISbTfv0v
2+cYbwXtbacpw8ydNcUfmX63D14yxwhXXoDkA9Bca0b6E2xfa/vVhEizixvUT3HpZlvWz3KTFNpM
eFqryTrdqx4MURqgWAP/m+mhevLZVCduCPvj1C6BPS6T7Y/OOMkDC1Xg1/0IQEMMGwxdPYCTUl1g
pzxdf5HUQNTNgL3uvYGj2/t5HgJm0GpVeZ6PZMClV/eONc1ibUkKH7HJhPyUW9QwF92yGjAM6mCp
npTUKDWr6FkYulIcXsRwYE5s3bfkqwDJ1QfhqTfRuwq74LexrAfLxpy0dexBApjKa7zg2Z6GclbY
mzjhYuBsbL18swzAaGsR/55EtsoUG8cTLbBGyvQ7RqhPECDoR4eLKRfIVYulPtXOdD0UlnrQ5P4C
ZS1Tgs2V3ebJsmWDN1JTJ8NE6BwpAUMMLsbboTZkSvN/CttjnIQJGghQoobaPds/vRqbHuGm4UTM
osyPWND/fAEQADlCds5JvFQqR21C/9JHhaENmUZ0URmzrIx6i9O6fBYDsSCuIBJyMMYM3JMk3+Si
Bcov+qEicq8l9bpDyeIEOWP1f2zg9q6oPxuYHE++h6w9aDbA7OA7fA4klknJog7kWVp8UivfOVAH
fehB/yD9Z1L1OWdoLib3lNuDzmedMdniLViyNmX9kUWmoNSpljt4W6wgcdsqCAUQujINWgVoCdDt
zq0ciMkcQV+DVqmYx4Sl2ksIE3fGMyq1BXoMcclV/So5T2mbiG2RZ4HVh3Qw6EZ1ygIV6dbJpS8l
Eosz+43TKuE/trnIWqzXRKg7Oux3DA49y3kTEyOt8e33TzF08T+kF7/nGif8zye/K7CQ+FxjoTP/
nd6CZmaYc6pHr+YcMNOEProO2ZhmjKs0ISWncxu92druOiAzKqVGPl0CP0tF/XBapbtepUaHH0B/
8DUZ/d/NspHRB43sGQPwXHvfrxVdeNMY6qzb62uxGIx+e/8MeU/d506T+FNlUTpK66k9uUDd4Q/o
O/PGePRZZdUPRqEn3s1yWjyLuLPZswZZp+eU4E2wU2GO9m7o+9XSOC/Q/bCOTb10yMrLZRDSJ+rS
WVjyX7Qin7U33qRk+n35jQW61jxn28tFHhdu9K5qggB1a8iI6XQLVvaikxroFxjBdsk4VBVIioNi
FRRhIEhtJf/rz49nBSA/ohE7NcrUFAtCk91CJj0L3Y/WvwdpiiRKSJnP7X2vJ6gD/UzrI5dvf8D2
xIXuo/c83FRAZdpmfsvTb2I1g1LoJ7IRb1mAAgDLlIRiNm1F4pnX2PEuinJ+RDloWphwncaLeSa7
uZNo5if92GS+CdBEC3dOnUdVtIC8pO+T9dDMBKs1oeFi8xwqhYp8/sVRXSLlnsxUcJdWW6HvkZ5C
ey7icQNstk4veeoo04oS29+0UWWio9C+uHErolgKZgtY/pjSHLgt3tObIyfva9RwZFwesZ3FspTG
7lger4r9X0sYu7YfCxrw6XUgtBYz3w5OG4x9nPrdmhr3nWyttMoBHIMdIaRjBe/pBrcf8EidmoYX
CUmPW1EgUXHLToruEhb2Zs4U9DZtAA8lWiQzfqIwAqHXP4EVD6p6ONYx/8s+mhhe7mose1zNToMw
XFUKWkQrPYvlwxrmQmUwEjcjoL84qRkCf/FwMI2ELNDaCTM9Zx6I0VeVuw2zMwBaBhP1gnWbUmE6
IGlJICX/SFSMHn2SaK1ykHHUJWniz0b87bJYl6tBMFKxod2UyEKTj0TTehoXJyP7oodJiKd4qaId
ktifOZ2LE8XOACf4IRTVxN79ZNe0NL69YhIvSl69AGQyGoWKTD80zA8ClfWBMNHilcKfTjmbUDSm
JN2YANjjkwipTfmxNdkLTeKJa2sqcdhVBhfNGb1oCjNR52UWJOX72nYZL2nek9cifcrcJAVmADms
mNw9OKvK1PqY9AhGK3p4ltrWteklNul61V7VSr9/9R7zuXI31c8iFP/3ohp5vk+qM0nUMvB0IQTo
ng7QiQBe26YzsnhPrC5HvQskWLPEp65yQx5bUtVsUFlg4Us15eUzfgYVIoCcy9+jJ/pQU+S/9huc
Upd0iTrjSWUD/CZ8l9WwiG+4mXHXd9eIrdlEru0zvco7qfy5XQ21zfP7ZdIT1XFMCdoRlkymEfM6
hNvsaAJxvyMDa8IOo/C51NsNFnIqah8axDy8+YzmUKtYxEO17mTxdDRDGK/KGEabzOKqdYxSKglK
hUvdf6wD6lVygJ8iEXjpJD7XwqBjqOXgCwNYK2LzlroHp4PKs2l4bXvm80WNORhF/4d9hnocc6c/
Gjo0erPtdpMMwJrwiMWxvvUW02/G6JhrdkWEoFvAnjQ7dEeS8LecXdDyHfklY3Czn6mx1tcxquXq
jJHqRQCo0t+VOPrXCcBHf6xILtlU1+JUTBgBgdmY5k532T9zOWKQItBTnojK4uPvmY6OGk/CACzX
e3zC7ShSVpt4wO5ubKpk4Z5KA9T1EmhhN3KbzdVsl1e/uFZoF9+HNPpjKLgl/f2CeGmSmDnhu8GZ
jV3pgmGJjeGknRYCBo6YN09uBEY04kDJnM37dYNzJYqroGAWXhYSkV6H4tCPoUkijXO7WtagQFGU
klRdVJwEzWy2UzHu8yDph0FDS+zbpfPzk+EQzw6iDVAn7M6Q/nTri1qAAtnfN2o1AFxpPiRl41WR
InvwkeXHdR46P1kIWKXoGt3bUQYI2gKLkWFt4dzUOSFUhAUy5mIxOxHK6gx+KrZuJRBm+RCx2E/B
wmZmvmgBzTEA1qSpAqP0rTqNE+EK/ktntGXNkH5YPiUXwZsmB+i7MZ31H9FsCB6q6naNKAVBDuhN
lpFarRn4/uXc3C3N0LoUsZubE2G4QBE1r7aqEvdbCUC410lRvnVaBNPGMZiebt29jzqMQ8TX+i+l
UOdwxLN3PpWKqONTGHojgeZOKbpv5oynZXRF4KRYO9gPABMKDSdCYBQlF2pnaM4WCtbLzX/n+4eg
NZdeHqBk1LYNbuLXVIvESsm0M0iw7dUATkbDBvAGVp5sFjnE5YFEJE3kJCEs6A5icykSdFNeue39
Y8O5CTlbCDTG8cj+2sADEi1KwNRqtinmamhQRFFf7IH4StAzN3lbPqeK8jTIOtB/4QPLpto7HLuX
m41L66MxMSDhe1oY1jJEYmu0c4CmqQOKWmkQeDcGMOFPa0jVycamMoZzOArIukhHTGnTm26UovRL
RjeNZPhQcfInx8aRcxdNYcapx0cdkA1Gk/OCApa/DwfX9A7cFrw/n/RoCo35Fnz4Qo4GAqBDv8ek
bHtgTMLlAAeSggrP7UPFPpV77s8H79TtOjANGR3l12GWwkbfrkzOOJGeauj7FBYAU10Uiab9JbX/
FNTmV1bvo46N55VP/kbODrW5ZSPJYqzPHZJSHVcrbbLXdZPg1d86+TvPqDCfEKaWjOmG0ly8JVBO
0+S3WKL6gxG7YeabpnBG63H5w+/U352CQmQBoK8l8ST7L3KqwP6vFdNLfZLGIQlUNhcdYN2vGg3R
VPI6YxBexzNNl5qQzeZrW6w/Bccy/0gy7hdOXXHqPbnWJ5oxR1BUGJGRe0vV+PvNGf2V7Cv/N+Tf
wxxQ51aFspLID7xtxxoQVEET4JZz91fee68S1NnB8Hbfa5mVPiQhBAHEuWlZJSHFlq6ttH7Z7tng
3fd1jo+ADpN1Jf+q6WWxTbagVyCZrweJOoDHV9OikcSdKFUfMhSE2DE4SOWpDNGb5Kn0SSnwydA6
UvfpmeyWJE0Z6Hhsfo4Xu+0d6SVLdmhTc4fWnZf2iY152B6hjrpBFbX3TIEU7f7dGpg+rG4NF4dA
h94zCNip3+lxNShjsQDGKagS2mqwVtOqa7inFUJjU7yNU1kN6hRxyPliCoiuVSG50kp3CM6DA/BT
z0TXNXpne2WEpj8c4FxUZvs9m+6Eo59vEc0FDOKjvj9w76glBf0RxHbtFB+xNmlIrKv6BpTkeAn6
Zl1xSVp0ZQNdaIHg9CqEZk/V2InvsTiEahAHPAJjBYshlm3PCMgPOe0jOXbmCZ4rnrsccI0PJCZn
VFwyULZaPZKO5USUuedUkAACQUnsIq1GKX9YtWOx7y290BM/UaVjiRXv/WzZJtC/5Unm0CAC4TP+
TLGee0dKucfkV042d7EFrM0N2frZilTXs39qbPtDZkxQu3bdA8Gzp1PnuEUF/lSH/dvlGi/HNPnd
KRePwtJAwcJj9U8QMx+g//pE2YIcdoTogJpRyhEM72bqiMxVJjyarFros2YBzGCmv/t6wtVp3n+s
26JXqKqvte6s1Ax4gVMWu9OUI5bNmV7O+LM7cSw+b5pUUI3bjRQ07PvWNzMy5ixdI+dIsvW+Ehnv
UdYfki4EkY3FlqpHKtG9M7cEf+rOUEolyhYCs+DnNI+OUc61DAbs7VHJ/yagd+0WiGg9XSv3QInq
/K9uGuIDW5faz4B0IzoamUQzzoNPft703tElkc7T5OGOXwVroc+AIps9eycLHocSU1wptLJ9HG7C
dp5b8xMEj8cluJ0vY0m5evGygSNK49AwBdlp3oPTb/y1csc9w/ka+qb+/EFFJ8VB7MPtpx81dUe6
HONq12pcYkyrihzvwVJnOydBvtvglI4Q1yRiEIsc7LFsr3fy2PVI/cK2s4etUG6SKTRaGUW0JaWT
iSOooNkYkgYCoOaI/bxuQ7oE9Md2js5DO+xDJX540vlXN6g8oxGWYPrH9g3z9xJHdCbSIbv0qZgg
wWIiPcocEyjSGSYndQUxNrj2Sxd3FhBjAXogHUsdTCAs3p13fKxblb+xVQEiGHfYudJlRP0dpQuQ
Ms/PQfmVz0ngSP50fEuaLjnIiPY0OMFwGPUiVrgxPMXbgh0kMlyrx4z0UXZUXXqTeUbX6NBi3D4w
x74RY73oGI5VuCaDDq25eWEFIUMOkBMq5OiMXnrnEaxipQSXGSXUEkfXNp6VgA7MClQ4ECwzrrPa
Az1EVzrudgFAT4DChilPg6Lbtjq7ImUIsP/EzwpgCv2fPHmVnl279mrDTCeBWNuHYBUm6QQ4RkGU
+ILbp8B+/0d/4WehbkUPNNzSb2mKzDGmzsos3hvs6FECSdeB9XFKbQVAeFlun2NNy/wFsI1lAWH1
KuetIm0KIRTgqttu6SWG5wD68248gSqI0fW7kpYeDwpDsu1x6vDQ1hgpqJ5jtt3+NWufZcxScXrB
olvG3CbVUGiE4AB9hXT2jgN4qKk3B4p5uu96YJYEXM5b16TEeY+F3kNzqK8wdAwNljOIVT+yLYPW
ZsCNkPwPbIpsiQcKUIAXPVj2wz6iREJ4Fs49Dmu/fLA16G1w0JgKxlyYXcTV2XM2AjW4NOrciWJq
qY6EscNxGY8xa2FVwVhj6dN27IjQ9h5oybtR+2o2s6H7/mbMIzkG0mw3biaa+hqRevnRppIk8XK6
5nAykOZ3raZ11hMEG1L/krCKeRvuBa5NEPsFOXfS072APx5XL0lEzZ44YTv2DD0QgsteVlnNlk7E
6C0aTDsyBWNr8LJi4wVCQF/ZoapT++k294ytlLrku/UyIQTFN/WnkUqm/vof59HnkSAIL96sHyr7
jOF/udSFBeC7ZZgX1L/4R8lk0KdfCUkpOAvU47gIZph8bj5XnsCXWZYHvsLi5q2H+aqfT/vVx3IL
MLwL0OMIR+rWoAoZpEC7h2mrOGQwI/9cTBppYAp9bdH6aOK7OpkSNDcBRkhHVq1wv2m1b5ucX3Ww
i2CDPn494mqZQYabu56zRvlmCbZwCI5tq2Y8v9J4LRweJB/50SWRLeOttvMWcS6cR7jmQrbqcBZK
xn9cbNlLSt1aRyJEXJ0RfRU34pUuwmA8jfIEOTo1T1GgBIGQ7Mw2S+biFVRDQBJ9hHuyv9iBJJMJ
Gx1GnSXd+26CEQQmGog81oNejv7BvU9fMZlD6HLnetkwJMVILXI8IGyhg3Z2Zg5lJ/uEgBCBUokA
Ij2w+OBxClzudTjdl34FwcUM2jTOIJYodtm/dLay7itu4XjOyMRUbdCnFl/qLkbBUuvymOVBfQcb
15xPc9Iw4lzlJ9ND1leoTrrXzgrsjAkzm0dgD+neHFN5lftL0F4ytVcGBeBpW9CFoTnznK+N3xCR
taDSaBV4IVt2khQ/kGWBYU346iObx9iwF/I3k9GcV2ZKI3obRtUw50qzvDMD2Oqcgc6Hbs+ygN0X
vX5l3yBri+YWZ3UaikMDzPdGJFyaAcnUSTdBA1YMW9nAILeZrIHDdOpEa7OQPNlhzKaDkNUvj0L6
ngAsuI7C3uXc5Wg2r76gZZEuAcozXf0rhn2Y29n8NReRzJb6xgW3n8z8bRb9s1FNxKoZX7b/H2eh
OvZYSbIwTFvLmjCy/FIYcZVbalzP9E+TPugsUoZZsEJYfM/0GIYpAYxnmoH6fEw5Dnx9fl2FqsAo
f/ApwqPFKmq3wRQZGrt52Ta25OGlEUIKTEzDaVBe7kJIE8LHuOPBfIlZhTfZvRTcbZOLuI/z9Y52
nHdOD9Lyo1hrPfO+vSOunRv9YE3VN39PgLwZy1FRLBSQHX7e4WgvTAn7pwO6aEjYAkyC4j7ToRD9
Iej8Zwzh/f8YPzZWxGehATo2Os1PxHwWAAFlQCaSQpY2fhKh1OoTw+xWdM2Hh/1JGe2OV4Hajqs8
aXKP5q2jAAR39qE+1pQym3ifUJlamekVJ+EdSR30F5CuU6r8gK0wT68LxSkQXjoic52aJciw6SLn
1y9K7bBcf2W+h+I91nlxmAOkoInN9ipphlMvaX9IGIEOTdKFrVOujuts7obkbegCud74qPutehCw
DOP0I9A08yMs/dHhAyax1d+ASNMohNGAluOz8oYNGa6NXYtEmiyL+oG/K9vDHwWJOrMZdPJLgT6r
9UrLTMPpJiBoHpsxShQ/GL/t5z55M6Lov9f17YZ8KM/QCXra8StgdRDyQyQVpirjYMBXQzPOFU4b
NrjF8cO0A9pqXdekO6L9ptd5NXMMRkUIfj0A2zIacNGPXtMd3ZH0WCHg/d/+PGIRl8Bk8gU58cKe
olXZZvfagZAY/J+CCZZAxvywDzkiHiFwbBfefDDMNCDXD5VmwIpdPJ+UuoCBD/aomH7BqkN8Pls2
YAjPPk0kdja5rvINgNlIgmrL6AAno0Hd2PrhzYFGYGg1bGql1p7dEHi1ZUfwM6TmjCDgaeO0kwfE
ivMYrE+rcgYGyfW4pbcgBMeoq0B8bXU60tdxizlh6Pc7uH4UOOhIqy8bL4gOCIjCVDrlmQvnnJnC
GICQfs17R/+r7dxb4qRGfBkVnS5OOMZpNAko5sHWzJetCg8Bv0eDdgLZUZtXHGh+tDr14gZCj/Wc
4mcPwWewDJF4BC2uSn9PPg3NZySzrh3+9R8yv7w9YcbIQ0+TJfJO9rDfUrskQqQTNVw3NPj9xr8i
8uLTsI2nV/0sE8q/a/1AyNbzN9/kH98HPQrm3CoQUIWOH9WDNnKNKmtGlxoMEu7Ob+df9/b7gP31
gKYVs0dR3BkRNuds+f1CBz89KHaw/gpaxOnkLlMDb5nj3cP9jJYFmuBbKQANLhNy/5DxjJkOQAi2
0HMBdE0rRWOe3l2ecbIi/lI4nbCVg2a7gnjmC6Zv/e0fZtpi98PBujvoUUTCoGpkmFRJrTBYQg6A
2A2+Vjn9PeATlNzuN1ouV3tpS9fmo5aupvb+xYAsMhIL+S8SlYKPww+9itScqSMFqj605v7ecDxs
8TwKDYN6er+AidjNiP5b7pLahO1IXvYXBl/M1K1F5FJISJMsSvScbmAL2cZafeNuUnfpoVV6JKRc
qyEBMRzgPVRySv9Bq4VRioIVbVJyB1Rq9+3TEYCgXP1rAByz1q5xEhTOddP/aT7IQnnALIZTjc0F
czUPOvf7KEmDWcRB/6O+/VLqdQcTNqzzqIK3kOiE8sgEyNCZ5PDfG2qJPkesPYWuBRs0JXsB15QF
6NlQVXeoiZZ9zd5H9BsmxDt7ybHzL2T0vx+p916ybSTymQt3UJZbSSttCJW3kQvvXMeZQTWuiGDZ
gvO7+FQMOce7Dd6kHsKZZoUN3tQ9xJxztd+ADOr2DJt/RJFhnYNbNEmRsh+jgKWwUXY+2mYj+nvj
j7DxcDXDLyhKw0bRs9T7Top5rMLbrkXIyj2iSg2w+f9k2PenIUFa9U0jzEiPr4ue2o8d/2zucMAs
Q2HkfmK7EM8Q4s1O1+LwKykHvTxZJipC8iWytI6nMFJDyX/Dcq2MBc/31oJq47/JfJl6ZsVwAhNB
8ja4yERd1Gjrtj/PnsINHF374f/QxWb3N/RVBoyZ2DWJr0gzK/pePP7je+hEG5lJrScaDQi/RSQi
sseSFjf9Mq3vKSM5l17yPeL4mqfh9iDAxN5VVuTq+W9RbJXP5UCQ6JNCINY4oW1xUpQCTxfqeg8S
+uPSthh6ZD75Ff+eKJnqtF1G9bzcazkxRtTsW9J/2Bm7DU8/yRpV9qSsL8qP5cXKjCFLiryj4QIe
hqOLDWL3rTD4KjIJaJJm4p9fnfRV3m2R5d2KheLNZ5B5IpqqBFEKpK46bLO3kSOhAsbtAqgrrra4
EOn1lbOMPlSfuanWOLhyZDNyVBcfunBRDAoE+/6Hn0mobuCvAxR5cAAdcPV7/9JcCTEw4SP3Rzz6
k6o64cMbLDGmXIst23BuXn7ggntu5MxDuz5jD9Aeu5bA2eNxZ4sHECue/ZIi6A+1ToKiDZ/BWogN
5K8yR2p8apTqKQ5G9suuc4zYrn1tF0zgXgNKEoaSl+Y413aCZkNx1nUHTw4K22VYHje0U75ws+lb
qEHyWjlVEkzUrqLlo9JqaVCqQ0d/TVgt+kWdvgPzuykWjL/p5VWDfdc41I0tTjoMroDR2XluwcQ1
qYpFM/lJFkl31GBQ+6y5Mc4q7TpvAPO4Anz5E7H4DApRu1oa4GovMdjinp13PQ+8hqZeFxoOTWg+
kTdXS3G+pWvzxLN4gNR3UM2wzgzCXbNhvtBCxiuLbGYFpC/pPo8LFrb9JBF+NxARKglAC30r7HiD
+0hVEEcptkaYh1uDh1DVBrZBvFwpGWXvYHs5PGVCWL+mBBdD7kGgLznVj/hytdCVyKNd8wYg7n+g
Nd9N1UjmfM1x/nHBbZgG3T26xfeb6clhJcFecsWnvFnJ3Zpi6xwHMM6cmOA3czO8EcpfdinNGf8H
RJPNb+BI3QtTcYDcqdXpvAnSRJ0ExvwbF6FMcKDlLpZy5Py+XNuqxrh600a+MKZZY2L03h6rz7Ix
fwfK6t5wmChWY0QSwTz4w25qesiaUSZ0Y9FGapvoMLfNIEQvmP4sszK0j25s53FJaoUtlepCuQ74
fZamHe7pVxZEym3pA2y5e/ozvKw8e7ahxJf4xX3/T5Pob9DcZUcAkb3nzC+yO28l9Y+2BxK9bxAb
InayZmvVFSTRNCKStL1xeaa/WoTxDIYyAFKZ+EgoL77seRYTVbsxdbqpLsh6MoszGVatsCyb/f12
b1zlaRUv6AjQjVrJ+f2/s9whgks1Xhr9FglXzp7Ib5iQrooxsPln+E0LFeN/kj7bU8gmTGKF3Mm8
13XhRZd5dAMlOHgeMiP3xpi21xmTnqXyt6feotqON4zZuwFkPL1GmNxLoq4f2b3lAoLeQOVE6P3O
Y+gLwT70VUp966gcaV9Y4eJTwWScYhGdnn+HsId2B/wVr2Sd9S0+jPSQeDGqpVsgXJ3+RAgPMf72
6+HbhsPKjx0A4cIqNlR+8cU2+euCH7/fCgJldo6OhotKMj7s4bbi1Hvgn4CvU6vlK87nWtikqKwZ
CBnCG9BBHTX8Fr7cLTdp91a6MZ0QDoK/OCyMbjQ+Sk3NEz4DDKHWtwlLwVGVqIM72xnarZXz9+z5
4oqdozSvP8oNnF6xEk1nFR7BgYvMpEKf6N4TboZdPRa2Mnh2LEi2J1tYYfiAx7q5gVRAPXNfblui
s5KRodjGMvirV1xqTqfH8rLFXG8M/Hr7BON7tmfT4qS9m/mimFSxMV8TCzhj375+CEeksSp/EYPo
ZJWx+FqhfLX28CIKXEUtK8mx354ndyNmC+D6Vm56RlsZv4bar94pV6PhIqzCdg6lDhN2TJx++VgD
WqxpEPd4mF1wLxIqJEQckaR6ZNBqsAK66tgRGbVGp+/2eWmyJHhv7gZPSccTN4EMKdxHFzPEJvfJ
LSHkTJ9Y+JWY9lasLkbh03HfXateIe5RZ5TnjoRnab6oiIYO0osJv4t70tj/AiQnAnSMw5diVeRn
pQlSTdyqcON0YOeoPolLYZcyDezVmQMwTKxUlrrMXJ5e9YsJF1aHCiKijI4Iy77bacEm0jfrKzTi
OG/rVmJHcUJxxBxtYHZFcn4X0mMZnogHcIvG4/SdRsvAjRgQQkNKYO3QftiCaNiAEMCuz48NYaUy
wxUGmPIVp6DgDIwT/p7XuNmA3bIbccYt15EnqHWpY4QaOELrM4JMIiekeDKi8l5YF2tbFWEW5AdE
wiHHAsXBVIGoB8PUm9sfEMLIEqOYZlxNtNN4w/DFm6EL91I/WJErGe3v8Kz4nJLVpTqHgpxgQ4DV
Cs22pfRLBHtsuePTgs2uiR5XxxtNdK+ldrBMAjq5x2s+kd8VUFTDFV402vg+lpH/12sfbOuEXnWM
Ogi6oU14UNeW7pXbTYoc5IIbd6NrnlMxqHmD0/ezXFMsvcDKYG+3Aqon15xYd9EFkEMj8fdocowM
IFqL/F/Xzh0rL87Dk0FaoIwIcXj81Qx8EPYX74REK2E4IYw4TBiy97V4IYVS9Z4q+le9EFaSAPLf
mnMKmnbiy+rwEeC7LuqevRissiwkG98k2dVEIuqoe+/aYpFDLjB+xerHnyMxkth+GE+FghEZRg5n
JnNZzphUHCR5gaZ82RIZHLb9P+fZgKIuAief8xrzvhC0VZ5BaiCRv59ZeZwma8olvG8d8maia9EA
1/tznRPTIjDP7iKrlYkMK6oaP7eruTUBVBiTqraQxpUMbk8atk4U/5CKwmqZNVBDVAzSednBbn7c
EtfY6v2Oy4n8eUAg9NK77Qs8+04qAJvM22hVU6jaW41DT9UEj2Q2ZW7bCKC76ZHds0Xt8lEtpOmp
hPrH3GDYDbqqrtFMb86twa85msZeZZzMGMTUXng/EAD89PuK4IPKEW9cEaM9ZpU/nDp8PrfJVgM3
Mc7SGdT0d8lucuW7SELJRKBwG47Q/1JLeFSl2uvUHJv8Tx4b5PMNmvjOLSl5drUNeji/uGme5KkZ
rOC6o0tdON6Pm+9X1dVut1ICvaSlLE67x1/lI47y7f51f158kHieCpLy0Rp+LI59W/0rTlgPPXyu
y1K2kFcowUOjtlouQK0xWPN6kiK38SpocpFd7IjNNXE584Fea9gZD0WGZmbYur66UDvIjQWbgEZd
P7987jbXvqCojBnTgf2EvA0LX5Qbqhrc1dbOCDAbhQykoo23+fjcN7WVJPw8qY+EkZBBT2TuA17M
ILNB+h0oV92sCEjwf1qv3YLAH1Gmw1wK9I9qnfPFzBF8nAKPK+TW7j5Tryi7dZw2gApJ6GjgJNWQ
oP20oR84yUsIB6MJRwTpkRwq7E4bSCr+pk8yMO5UkB3INJsMPFj7l2iZZyvggk83hdNOeqn7lwrd
lS/8x42TojSPhT5cmA32a4ZOKz3Y0NWnpZu0JarUL9TZw2eaOlnu780VQzvWP2a/+R8yqs9hc2Gr
h6ajeLmo0ifF/LpgT8w3yGn6OHjyJLSUlKhU07cAHG+d3vD9NdIjU7YHQSuvHEeDf2edFeJ2bs94
CMPbtDiDMyeodoKQVwpFd5XmWNht3OOy/dS+KMopv3OBTElqRNo5WrO0WbKgsKf2jZf6Xeiy1FC6
D1hPzzT05xLEVaoBra51k2fUDGtvQAuX7obvLAKNDWLsl1g+q0rszaXljz3MZu4++9oWH3bhlI9/
4FmJHG3MhefYiXy8/fpfWDQcaKoAls7s1quK9wyVbYiF5MiJBnbNkau2jRgmbq3BfXv8zJMFlZdl
d6oreHLPrylPogzku9XL2dMJ100MefZaqv1CRTrQ4OoEOtgEbpW1lveMFGUrpfqdwEbcG/7qFEhU
IKXShvuVmlA75j70c9gCMsvwaZzoKBySM2+Sdnmcg91DLBs+e+QdQhGgN/AQ9cMwQw4t5pd4s6Dh
NR/WTN5pOgoWQ6H+yFS7w3GxIdhQ2Bh2Ir4gQTOtLRKuwRkMPs50sP4iO1CFDqO0AaZfWCPgfOhY
Dgy7MgChVEfa65BZXzyK//h2k+NVW/v1F9DvyhB46VBEwD9gMRGIBH7r6moaG9U6ygYCQTautpHg
S7dmrzfUUKV/RrHndbZj5C2MccmSnr4x2FLuqcoXzaCzOTOKBPp6s9PiJ5TmAPJ8gTvHZLEmD2oO
iDvTWoVpdWcFIRR/s9MyyF4vccLq3MLTnIiqpNQnEKuKI6bF17vM2V4QcmM7iv3kt5Z1cEM8Fi1c
3ywifGsNoQOCi/0vNJ8dzc9KowH7awWHkQ/mM9xMJRmQ7Bo232S4fTdIOswENkeWSQCHjS6XJnJx
+bK+LpesKN4K9s56E8liICBvHqRxK+heOqixvjRtHHJHwqZEGJ/Z+4x1OpmhxXouzYhnLX+o0Nqv
U6aU6LxGv6sQ54Wh47bmgc62Lemx3K/4Txw4Wl5snA/4QTRVcd7fKzI2F79k7Ex7hGtp9HYOzs66
3CjUNflFYIdonSJJ1WChBkMr5WVfO82Kb5X4LeEH5Yc4B2M0rHXf2s5JGisOweYnGyGGFqAAduV4
7vatCG2ZZwMyAyDQkIgLpfrERWIf969jLb6H+93ZPV+GkiwjJT2uZk34KtQMpgU5NSbbvqkwDHyD
hWgXKM94U+Q4QdofdmSTfDO1Br9rn/2szgC+jBjtRXrd7cLdCLk3B0D60Tes6Tt9R9wRWkn4XFKS
kx0tiBaUcaXiHp62YhpvkyjKzx3b+SeR5nDP9VokTUHSHSVZ2FTN5zWY9OYIQjK/bYezp5pvBqPT
3atZzeAqUIttWVmHwU+sZ4MlEglocqWEMxTLhfytHyVxKvS05/1Tg1qncRJOoJry1XLLiMMe4YBO
jDBzZGKhMPcDb8rkP8N2+mbPlVNMP7xOvblNXcpcyGZyu15IV3wRH6G7JHpL9s/uuPGNlJHK8fRS
/bDKBQKVw9CmTIIjSXiFMZZNRdkczcpC3VnAFi9sc5YgYK6rP/JsI4iCswZKWaHlvldjzT5+b8P4
9xLUIEYsn33N/ZOXMS7RhFfB2BWuANzjUBl/UAdkaKCZxiI/OfCLDzxmkV/jDBnO3D69Mo/XpOzs
3WmLdOfSeE8BB2WVWEbqbkeq0RJhJex1VLb8WZ+FNxrRVPgHYGOXFZkmfk4XLAcWwmitaYq23Cc0
uF0mL5BAXGdyUPEzNV95aSmZn3GIxpDAEV9GutoKhuo5keRJC9BBTiwHo6U/dptaGA+i/knkxxnX
N18Lec9QKJDhESMwZQqYnDQW7ehem6cOc5yHaZA1T/59ULohpyVRzbEvgxPs1kVuMgplGXMl8EHl
+Vkpk1FTaNlCdD8wbeYFXKF/eFf1LyvpwWLdJcT2gqJgF0HdOELee4/1l7tHsjRifNWHIa5RAAtz
UpuHFgq+SuOExY7QvsSEZWyJ93KWgzb6Li46nz0zxuvn66Zw/OzUlF8Xdu2l2KpMcyfYTTtewIr1
EFC8aXt8XIIZc7VO9rQjjUzvkvbXUhLtrJ4pZqAXuZoU2W4mSDVmFHQ0tnzKI6LgzPBjaHwMIBF0
1Gkh0+PQL1RS0ztQGx4WwczpvjVjKlSJ4WoLoQ1PD7zhP0ZpeGc94QN9wv1rV6YsQM/9GavGga4V
0tg2Y5aN5C99vPAppML+kagtB4915HWS0tzG6yFb4TPDAIK+Ie4GAaj17lilTlbKlRHbKstUPiid
halDQKoO0PTY5CK+BAaQ+fCNolvPEK4KeBwWgFa0NAlGj/mNurhViXraUSoeSZwiRu2UqrgPBZiK
s0DPyrUMmqcru83+eo8oMrEkw7jw3oPiA6cwY3ScqIHLYMVHveKlU4SqzWVxZAIy3r8N14YYe1Ej
mVaIMiJ+1rkeFrQvUsMw9edSi2jaL8G/qHmxU26XeExh97yCz2EGT+kjJAbWH/HVvaMu24hKjx28
6chTDXBferDddqXKjG0XQpIaCpRCW6T9pZp/j1cHdhZVSpbJnW/rIJz5QTarye++qYX+rblfFUFf
1WseFlmdwf5Li4SWNlj9IC4H0fA+WYUp5p/GbSIjLlsEHI4nb5B6hej64UuQ4bJ8j6zAphUrMoOO
EgYn82BDeJqi8VDu0GIRKmSfv3xJK2XeQxf8kgUMn00/ZiEmC366drpc5xQwaswBBwEGKd7dCfHW
/9uDua03TGz4xX2CuhViaaAZBC4N6fkBKYE8Hw4z11QNfi9MwUAIzd9R31w5Q6FYKaltTTkp80/w
ERuLs9wQQgDoaX8eknZdk/jWNmfhKkylhSLfFGe5RKErcoZvi9yMjXHd5UBeYfAo7B1zGj0TgkjL
nm8wKaYZXZDSiWVI0dHbIgBZ6n4Hbk/rNiStLW6utlBUeIW5oKOXxuEACwZBrKWH/Fj3iuo4YZX2
nxBe2VTMokHMI61mkbGbhXorl8gqgOSglLo2HzL7kgCPvBydo2wMoqgC7efozjFCaufunYNsmTWJ
xR+1J/I04NX9wzTYDme/g2cS2MC7vhSnqiILNwBAhKFTYQk4dRt8MeRaTWCDTtA/sDVU/cgddqJB
CeZYC2YHiajoufV/u7d5h5WINi78zUWeX43lMWPuJJFM5OjpyZXbGbRx+YD9c1201yrmJ23UJy76
a0+L1bLZ65lgiVVudTr+mPjT008t8efsQdjJ9lOGWhyMPZAefb5h0Or7zAvhOosCXL64/tcT3h50
LWQ4Uidt98HlvTCLnSpA4ZnbRRkmaSiEEc7sUtyJYPFDZul+0w0Qtejv1L/rmAsD8SLjA69lmMbe
akPNnCJMWxskRsZvj5LVvOQ7q/UYmiBTIv0pHz9jTOrVKikEqSzxa1+u5dSof1AwJawdqva8lLL8
BUWXCJ7d10WPgeBDuQ5m92tRibK+fbriEYTt5rOcVTneFGTwXTK851uThUaEnZ9Dkb06zGQ8fVsk
SLBYFYEm3nMaXvWgzXGAB9sjOpyPneXH1ssGmpywhKjGAxvRzYVhl8SKZ3q4PRSkEvs6KfyqzVc0
/MdlNczOHgKVuOAWm1VpYRtLOl1xLO5Y5J/18UkNDOX9FDlZBnqE4CtgS7FgSC3t3kutppaH3t9P
puFwJIUlCiB8dPW4tSkN10hIiJQc3FRBy4HQRqs5O2TWC7zGeG0pt3PJnPOwPlFzsPG9L2fM4W67
kHlYwUO7ApbrCv+BawjLtEWK7wyAE9gvkQbh67HhUuQNxOuYA/WJ6AyF2ebaohFvcTar/DFls9yI
9hgRM0MhN7WQ9Y8iV0eFMCPVGm89T4TiYGgFgdrhO+FZe2IvoH9CcvtrAuqXOUUFmuJq1DUZXc0J
n4V35wy35JNu9FxIqAMTlD/gFNr9DmwMO4eXGRFiMDjxdG+1fmrDCbIHy0CDvhN+Zop8r+Nj4ELy
xZn8BV1/0bJi8eWfwgjL39XSF6zDceV/usR4nMWnq0a0YqWZ3A5+W3VR9KC1fU3SCiliVdzkE660
yFZFQwVo0hjPHQA2pFIhhUbM3QXqOXEh8DE0iQyppMwXHRPW4C2RiCa/Ini1eaNxofsMWbwNd8Ex
g41zimaLsQ71Y7BogffipgJ2HxhWaeGXJrP2MqloWRUJRABgC4KVVmBGBnsJBZCi5H78+PKCbeAs
Sdws+z1OXn+N3HnVsYBD/stxM8QOcBQMZDH3UUo/1BPZTkVUYb1T5nEjONf/aHooLtVNXWTdWlKf
+1/w/ODgmEVOS4UD26/IjrWYjWNtK7IjJP8c+HjiKdSA1ya/98Vgrjw9O/bBXRlPtNW/qlNbP/cX
NBpBzQKInHlktfUNiCnC4AtQnrinD+Y/EH2N1HhnkvscpsadmIyFRSn90H1fWg5w/gpX+5C1zrGy
c/uTQhtzD0gNnSsJqU53PldG9fwMgMSuNicDhkIa+7eo2DlJusMxWCT1DqjETft+LB5N8SpRVGLO
o4geuhK65mdfTrw4jCC5QOkeUExq3EAH9Hy5Sf3/3t1+a42CYs8g5EEHIkBQnS8kgmMwgL0hZRRm
kP4sLRBe8l874PqXOjySHrP8taiKtAeV0ukQlEpm/6MoFQEl08wnodPTb6WGsZccPN0FfoZKjGNC
+O2/MY9gaJfbNx9SyKlzJfJLsLHiWw9NLT8fim0WmRIz2dOPbZ58vjBXqcU2sHuthse+tcil0dj4
2kOlZCimenYTobm4NWu6oE61EQ9U2c4EXm/kWAvhexsDosTCcBH2MOlZCu4JzHZC4CsZEwO+yPyc
yPnq+LvJP6mn+PuGiLMpiDSb7mHel4fOpDCQs0VKAheX2ceM0CBxrTbTTIZu65VpcFp2F7JywRXL
fAdmUj0QkTtuDGlVcc0r4e/P7RxLfHeRbogN1ZgVN0WOFC8rn4pHMWcKk8EPbk8F3FACgt8fMj/p
ha8v+ROOY6Em+kltYCijQFHtcDUsQxWCBOoZOXOTDUJXPMD2UwJtZsocGmzHgsT/xXs1ztFOHx3O
SMLwcRJh9NLjOt/p0ZqlPAc5xS8GbOfUwsYDbPObbF6LFpobJG7BmIndk2UNVb3h5SgPgYsUO+8J
8YUICLwMZxhFftL5yxMWm72AlF9RIDT/dd4TRkpIOowDE4+0Hh56Ld/EOyKXpNSWh8KA08wUepdY
Ye4S0SCACuyooFI+tJWlGZEVIfxcLp7Y7bPxO4HijI2lWO2Qr53oICNVjw4EY0/61KYYEhaBtLXF
7t8NSVhkGf3h3NdX/OZpEEK2xWAAtLdwJE/z9TIS/mccSnnOuqTprejbXvhEVwqU4/qNm5U9Fg1r
HTNsHV2hkHll/6t4tDOc85X3oAZm8sA3W8JofJ8GUt4/hVJ4bkm2SCF3Q3xrJ8+YYCJDql3wlF6d
XzbkZciHpSVwE9BmN0zMQoubtNwDUm339Cvz3Zn4aQJz/zmGejGLrYSzSphGyqyQcTPmf6YAKjtX
VQueieWXv06LmJNtteLFoSaKDPfvDK64WVo7aFI3EyNSJk/QMmfkqaM87ccsN7V2GNbbkGakj9pj
e33+EoqIlnZ9MQnbCcv8uqGmletbRZJu9tfPJPRQ+vY6FcgnMODWH+be2/8IzNrpL7IPz35/gE2y
vjua5cPPxGKS9vQq6yJkTcKeyZvtuu943wQiSr4XcyGGdvnnEDyB1QOxMAtC73ZodckxQm8pqVgw
AKvWZVHT1HhlftScKjWPxQSKtCjnaAgjV3hZAsOBV/271bnM6LBGpaOe7noGYyuSM+6SEbN3FJNp
9H1+Ipp47jJNkjX3RPM63kntBo6pbHjJ86+1PHBeeUMWpoWaIS5m5wp9K4TlHmCknh2Z37IZulDa
IgCHWvI79qIVKzhYSWuHToxyKFZIB7c78EWl2rDLFFMZ09lXITRnB3ybLFFomlqEuAQ8LczM8D6m
S87972HWUWbNxuG0YFBwJl3rEygr9w2LW6CCN1wyR2OY005mjPXAr/m3PzQ2k30NfaiX4rVElcRG
Qx2J9T9P9vex7v86/rC92+5nZSK+oBRO9caF0pCZS0IMPtAHS2MVfs+78X3GufxFifASFqm0jBnv
OzvwaSxgJISU92go6aQibSWM2zWcMDv/BWtYg1KQ9ur6Ej25e+eWqxfiqu8Qq+HrhFZSV4olOKUg
qF/chuOXf63UdmYyg+qt6AxTK96rqjoJIfoF+YUMFHCiv/iGcBNzyknMqBDT/cYI6Lx+djv1aWF0
Zqo5loTy3464mtsNgvVk6rNRCEHaEFaEysLWksd+8mWzzl+y1haYboBToOYnuTOd34Wge6g7CK1P
QbRn/Gz0kdhrynQlnvFSmwZmJrvTebldHwpPGxpwaqzNwXrJdJqRs5lLPL0asgh2FZZjf9E3vMW6
BAKuSQBkw+v7GCshuxEszfZD9aWg9kCFMw5zmRmQHy7cVXYXW8qWkVQHdBmQprUvLUBnpGuPahaY
7uY7c3Gccgz7Lj8THYMqMZu4Xpt5d3kt3EjLvVRKbuxH2v6Z6xrVBePM9tfzFhBV3aNjJZCciMgI
PDiDdMSNi6T5pT+ui1xUo8Wn8YrymWYlKLNFDEmSyxgOegGIN9kqIqPU6VDJWXaWTlNuKh8H+Ef7
HfY5N5+JZSdsaFYBXbl/vXje4KBVISJC+Qv0QI7QtxGXzjdH5NTs0VwUFcpmr5VVKng01BZ+oL4p
wgTcQvqgrSYYZ4dfmjmG/OLOH634o9Y/Ih7JNjGQ3mEXVnFldxKAkD30VW6he/z9s730ReG8uH31
F7LpKo5KDitrx//B0Mi3e78dzd57PUtJVAGBKyvybIVNywAwZcolJDXTSLcnIJHp43z8bqExlS3b
xvi72i8ezbItkQyOSZmf288HZE8oCZt4PwMaLvNCS8oHnYlU2/a84u+Yhg2U5oP8v7PEosuMozrB
rhQLph9PbprHHxU2zzP2p2rW7R1wUZuD3omrsrG5w8gwBCtECzhTe8OA7uW9cLjtgNlt4H2mviaK
TrPGSt+WDmwig795E6dv6y7jYYJBljtS/IikLt3J5JZ/UdO9InAARcBhQM4sYGRFeTprTf4D15q2
N/XSJw9gBmtwWo7ULk3whPafjpl/rU8ay6/iSeDsAyC+xnbYSmiQf/T70SNz128eeCS4GoCYTDhc
5rtZmNDXWXIZaqejohhGqn29iY920xeC1euSTMDyeqs1ylsggkr9q5ZKM88GtsqRnw/neWwUv/wA
OVNS8CUFvdKnvwZEnVYFRfRFz+1lsufZJbyfym/K+yAT7DPvUyMIiOsPDfyxwBCRjiUi45bsfeb9
AqU8PAyEzfqZ3qXBPwcXwG2AC+3GuAQYCZqEFfVnfU29kpFOAFtAZ28Hek47PLclxS0wPz/R9arH
tBNwWvS2/4VV7A3/BGCvgLtpGZmoer0mBR1/gwTIGXDw6OaWpgNuYkLOdciKMGJcyzNHtk+rARjL
V+C0bLdCOtQzvjAfLKBfCv6VniUyYQx+GhEJGTWB2j4siUa+wAP9cP7AjAeTOiSuwqnhPR8W48wy
Wv+3meRT8VxySsLWAZ0/YhtGV2AQD3me4kyFiRWS+D+DWuCE/ozmueILakUesh7FmqOTyHoD0FnG
oUsyLW39EYgiAtsWxUzP5uxLPpQys4JX20X7ZydW+9wKgbKNs+/RftiYcM+XaXpVs5cQpFk18YrP
ymYv6qzP7wf426rkEA2d6Ap9VkDi/ZH7iX9EFkfSaQOrncayBOxzPRxbWyu/Ty/wyFmCG1266BJ6
RjWXgEAZ5Gi0sLTWJYblgknBBZAPMULfzCStHW4bzRZQyPbaHj7zmp2K5YGVZhy5JhCb9kefADx+
65dv2OvHc6vMhzSj2pjbMEso/zdgaM3L1scAEEgCUSZgRBXQFar5bzSMzhIhoEosowrHB9FR88xv
qBpq9J/xai1YQ/4zzTxFo/lsWTJsXiPF2kXvW8bBor6gXklIte7JdpLwxKcqRBjT7yxNzAoOyx3i
TesBsrBaEcx999x+tjMK1gm6Vm3g8IW6zy7A32FMI+BU62wxsxMcGujlEJfYbZXK6xzcQp43fk5C
Y1O49yUVu2eNDox1Oy5RzC7E8uUtqd4hJWp1a6SVA7ZoHQ8zFeVrwe1IxBnzoZppIuaUI6U5flio
UbHKfteicySIzyw9F3O9ojVlyIzYf0veBtTzOkHcM+uzjPaDON7/J4Xl2MivY6f2KnlLsE2ztSIo
P5jVziAG5hpJIJcOoKA+9qp0SA9eJOvQN1EOEpeZgrB9b6U/ABl3j1Bol5r/CD+heVpIu4o7658P
exokOew8ZnBHTrwiYNuRoYz4nAod8QWsQrcYfTo6l9mBRPAk/hVJ67J5A6SNMQo4dH29tc/cWlMY
/ZivAcwnaPDYOIoAe3jCM3/klrjO64hpW+uIuOQRWc2I8OSMiSohAQJnYlBXY77CWPW19gcJaEqZ
D2uShrHNNzzDwuGilD8NIGOrJxj4xM7BrdNF4brull8VjCaTXfTsoP8OuxeG9Swxtn8Uf/Tw7WZA
OWY1p9rnKckwydagQqoo3HCSEjWkzEQPxLnAcX2SOi3Yk/niI4JU/IBTgKFvniOoTSzqYlPs/UNv
WS9WErL6tVEgOKi1oCm2vPlg7ouvkjDyOwMmoMRKq7IuEDHo30hIAePOZqCarwMdwTytbR8+157j
UPXAvuYTkTn2QJnRgjEicgx1jHd8NtJwIGFobt5o35Ib9579UJPpisACXbU0B+b2G60JTIHgsBqF
tWMtaN1WDX5ky2CzO0KyLDdr200FBTNguPPog+ESfxqHNsjByLOBmJWk9JvqXYJqbELWMzzfDVPA
1BAc1tgHOWZumqqVyDrbQ0Vf4yeKZE+jMgv86JHSAubijmh/lF2fnLL+Un/I8pxEfgGjz6knx/5q
Ee2NcOuETG65Mk8K+fJvlbaImUTwvufFthSM89p/pylqSOE/8N2/VekePUaCXrL1+fT9cDvsa3Px
bi04jw/RoRv1MAMAV7Ya4Hrmlo9qhGnaVSjxGL8q/PXQYrfd06YWlY88mKDXSP495Le2Ylk9kjmp
S855i/22NOsmjNIM8G5BqDOpvI3GGMG6pCYH4HQ1nVYIhvY6JuJSSCBLELkY6uoQwq85ZR3buMRN
OZvqeap7e/cvXpUZXmmTg5TAwqaL5lV8jZo/kC+JEXHiJPuGX1DOmR6VSXKZyHoS5GJdjKispQpO
jTjdNANmBbcsvO03ZCK7vzhY08W+Obn0E7e8bUg/zpWUAZQ+d+LENssTsfz+2L8IaMmmC1Rphy0Y
zJw8guLokHWkC72KiHban84ex4OORAt9z+Sc83VlMyzltclVicIb2B+55Q1Z0ea892Vhk2rN2WU+
UJuDkuvRa+PhQb8N6K82ghnffY2n/JB9Dt7OC0kN5u0Rh7YbSq7bS0xl/VaES3m9c+k5oEsttpHP
ES1/bPGB7EisrPs8pIeZvt7gxm3CymVgh5Nkn/p1zZgfqGRtCJC0wVY3tB8seQCS96xDAFfqR9OI
xdy4K2Xa1kYu1tqnYto4jaM+utckkRQ7emu5ivFHMiXgX7WvCm32TIJzRqjbpxT79Oz48VadYGLf
+0is/Vq2qIqGrssjVo+JxWBVdo8KpvY9otfeSZr95CgEyToBYsbp8Ze/Mr2OHOv+SiuWqy/5AVzi
762KaLSrOHkrUqfG5abbytOSAcFqSTsrAvzVcfjEdqk7xy/8FNbKS9EO7yZ3HuHSQpIWPRoqTi/x
8dXm8ACJnOs/Q26nPJZnYVHNrEtqF0Vq0m+XB7Hmr5Q5vyU06Iyg8oFnCILnRLChML2ifgdw0roI
LjjTv+yGR7D8aaePfeyfebQ1lR/lkA5KdUWD6M4mM/n8CgD2jOBq3kakcmu6ZD5GOMY2mjWQOYJs
Po/ZQxwUQdK5M3LfTs0MFCs4qUz7Y0BEDNvjqDUVaLVBNgKGL3jW+LVaNUPnu5SVdyW5IJuFyDnF
iZCiCmphoFtumQllwWPTc0VZ+CZxlHreoaCJVR+vaBObl3NHvVT1P7lKDuGxQBLVDebT23TBAh67
oLXuvfhxkIHtyA8AZq70sSjcTSCm+cddDcJcVSYfLjJ7fRMVtZdEaV46L+MRKnFp7nFXZuz1vORs
KRU0bAwWUhI5zdNrVePV9l3Yzeof99reuMnMkhl6SOeSnGIfZAMqc/fB9Uggv5e6xZEloOA7XvAy
+JjTEwviJvRWoT4tIUyGSDLOOS+G4mbsCQRBGt6/Qk4ULaXNI9QEQabt0CFuf3X2dNFm1U0dl8r3
UJIf/lsQGQ7txA9vIpWNM4Lhr7TK3fWQlRRowmy1hz+pLMecmx97wbKkEoemhLna7oaVNULESdDB
O5TCwG8njeOIK5EjtM99yRzci6Tcb6YVO23qG62q28XTrgPdhO5yMhzz5X+pLLQx8GUwmATwYHo+
FYSvXcONtkAsWGcZiCEinEwvl604REVONS6IHKYhN7/soY3J8NpjnaY5gi7kjIgSteuhcc3cVJdA
l0p2gBrVH1NkpdylBmqScW+pU5agynSYzQ+DUTNXIwtCE9Q8CL7LvwhuIc5VMPhzKRMD3BSluB5H
69ggCAYwu2sXRutdDNciXllZaqwmednD9ZGX3tIC2/V1AV32Sb/G7MERvgOzUdLssTc5cABZasbB
tM0ilosT6o6hUQKubZPIY6LjsOgNlRYjdAlrFZMuXERnKtRvennOZegA/iwMNN7mlxxhm2eMdpSI
VYOwQ3NFKfraSdNNSVD7hfFRJgNJQFs044Mdclu9QYbGq/ZGJA35rY3Yo0GgLaaYjNFm9YOA7Vnd
I1PffXunF7TE2O4aUTr581VgPTmHYF/DjrmsHkr1L39JvL1ZVbz4ItLO/SruTveNOxlxRAcIOhSB
mcqh4qg3+2VF28TI1Dz9z6Q10Q/WJHP+4QxKEkQ7SXcwDq+WLpg8UMfQez2Rc/WgSFq9Uw0C7Vfd
h3Kh17zh4cbuqr5z17nPpxE22DkRUAPLGCCFs+gGS2cXZm3JglkV0zErcfI7wLuegtMogpPQabDx
fvehVf6up3GxGOV2jiWDz8WTyoPn0A0ezfw42ci7CfNkL1YbxXadHmjxXuurApHW56G7LeZx8YOK
Tb6ocHXZq7jvhzy3vWSE4m8bFZkncj2vnQNRHmaZT74pLOq70GkuQBstrqWPZAM+whl7EFgwZJKK
rtEdSsTEbCj/wn3/lERScMPSN2WuRb0Z0nZc+PYUT/4SH8yE1MdYGCX8O6ak9yd+eoo1aRYMOWTo
DZ1sY/jWWwSeRYhbsjJ0Ilqal1Q2S35y3ErTGkEZtGkpe/kcw5Hs02QejF38QarzgWZnKUh43Hic
+W2QcGMbwMpLrnkspVZc7newgJ8DA27N8HTFtXS0+5UQoh546ohelFuQuUdUDudlg13c07rH8bW5
No/q65U3vZTqFyJ8Vad1tyBRDST6dyCvfbqJIhps1c3Z/yP3pOC+odfel40YVV44VvqeE7LsZ84c
sE5vExrs0QFTi83qytpvMct7fkqRUbq4HxIpww/owgSFxEQ1DmvxVTbBBV2/l98fYnWoqw6oTKZF
AnCsjc52zbyomfgqaW3IwccstIvh59VfSrhhpNsjtK7hsqqmICStJwLK0+66wr1AgvcXXi4AsYhJ
s8CfoZsHtufKWYsb/EvwSaBLnLpSiEUiczqMWwC9ye6/muw8RgZ9nc/8kvH4GbrDIhJh4r4p5H1D
qEDXSL913YLN0zMahYEszFGkQ7LR/oFqdd5hKpv+/jnARGY2R6xytOVQX4V3MHdPybxQ0vWHMR4M
Flhjw19yrIWP82xnjwxTxwp4wv4CpslX1AStTsIgBrt8puyIysj9pVV009GygiScNxAOMvIvpySq
iGXyD0KZWe8iRqKtgs2RUjLWj/UnhNjR6swtIqUF46U4aMZUNYkPJOIurj2AhUWsheqPyEDVn7lG
7e4pQFoPzc+fspxJvRZBCpLbo7a9vtgn+5Q7T7oK1ITqZxEs8dfiKJPRcumE4A/FTCrK76pK+mOR
dOmfIC/srwYraeS9KiC0Y07B4lS267/KOpsPPy5e2cKRssbg1xKwFN5KhgTEmUJArLOoxBDYSpKq
88cDS++Aqw8K7ORLFpGlxS4MBC7O8we7ShPK3PMjEFurjMoidwUFtPJbJ5bpouVrPfqKTMKkFEe1
aJuhf8WgJQUgtmeQAZx3U1UV24Cg18kJk91IbP2GBLu2QZlCkdfHzBahIb5T70UbDq4pdOwQn1LJ
xpk7vpcVmLXzPqE4eVgZV0i2JNcm7ED2+Ga9XTa7Psq0OrntU2XyWZAovcN4ADTrl2nD+IYl9aWV
DdYAQ7K8SyxEMX4NS6eLAnkUFHhWqbrmyTFPYnjbKftl0JFUFnP5ag7Qom0XCG9HjTYOP9F5BQeY
NFCBIqBDGMRhuf4AwU1koc1jMY5qxPq9cbhY3iNrD4LMCSmkKA/zXNSMbvjoxmppx7Vv0/7wZggL
18hCItkbY3yZgxB6iHQ2WZa2uxyDZN8lXaq2e7nMXZY5KQjwYgpj0gWlhIaAW0kMfsqgy/cmNuu3
VuGkVg8Ud9tteeNt107vMmc+Gn4xHwHt8AoysUFiOtGsD7U6orlzhUWWztZPB123Bb0f+X5MJ/XI
MZcD7ENAE+b6LXuoanovvBtgLdtkcSTtNxJLAs0xeE0B4mj7ZSbZP8LNm/jlEEoSiJYxUQ03teZh
R/ayeDoZSzkwFudmEuVYSChTSjlzBuV2sIVpQwoPHqZQLOcBwZYMqhnhusGlhIprQICWWRJKbwjU
ayw4c/g8suHSwO20Iw4c/kTgWqKpBp0cKYi3Dbc5fF61nkp97wlORRRv2dqV/3RvZF35XD2YYHai
wNjbVShQLpHb/m2KuIW9P4v8kA1UMzCjnueVNTxjgLfrnl/MW7N4HFUM/d/8aNaA9uiNmkaw67Ex
5Rsc72GDs2UEcQselDM+Cj7J5qDOyFYhDqhrgUsyoTIQQcQDV+Sv0mOKkASg69hvdk6shzqVjSF3
IpIlhdepbk8tzzX30bm2QLCUL/3+CDoqsa+NQHZ9xWSIwgMNGnFi5DES2GhKYZN1n71eKtCnCzKT
Wzt3J9mmU6eenkwMcBlVayYgJt7IUL4Pj2JIFYeBewG9xtbp+uUxvahAJZLt9BHVzRIOObp8HIfw
4rG479Ir+wRegnE3uoOUWraX/v/42+7lr9x4jLSTA4h7u04A2P8yZQcCAl6FRfEQRP5ujxsA/uQ6
UwbR2fFogbavyXk+1qa2Lw1SR138u9MH9gZ/Cu5BVpsAzSroCEkIPGRd3owk91usYQY3IDS0MBZp
bC00LVTgdEWT3MkPqONH20kuZWNRi1Ra/hkdy8y5+QoN/PDgV0bvpUujj9+qZKBaC2aGUSPbjEbE
YVvlIWs8vCEfdNrPeVICC50wJaOHfLZybsqMmYM1oCo03qqhPg3rtI9eACy1t+oF8w0JQUhLCoGs
JaAnL0Wb5alzLAAH7ZNmyjeyXO1sO+dhYOzGwYES2zbtyabJdaTHySSjZGREQt7Npf1H4Gi+YZJI
wKq3riCDJxjlues/p5iBk12rMiDMO0GRNrfJO4gUCwxlJcYKAAEVXsVTahHDyaXlW4/qNzB/iOJf
DO5HacFZqOKjwL5Xa7sR0awEWUgSlmFM/ZCai+cHt89x6OlkfBm7yeplWon/5Dm+zKlspAoDZoFS
UIhCaTm39GCDK2dCrAbrhmGrB/7uvsbEU/OrIxF9vBg1uBdq7qFa5jrRfX8nnMX/1nKLqHRkP2pq
kDeBE+qgJTOdI3Ew1gwOtWs04+UxmSnghBspEH1Ds5NaHHFvtSbFXXgzuUldcLu+t2oarwStrkfA
kQiWyD3ALcoUYn0ziRPQrVUL7fJcrzOGq/5N3RrnEDYj16kZ3jHIOCReNN87BAvrBuO+vokO2+17
CjH+kRgP+5IyFbntA7KjCAqfbR29TUwzKcAHG2V65tsFxwwMyWSKPtYS+hhvuN4/hXyfYPPjs9dl
UC9drvvIR/kN2RykspGvf0jynBX54ZS1tZVkTQwGhh18cb8dIp6JwX6zTgy/UMsj02LuymUiZVZi
eTd0s7X+AkB+Y13dlqYzWj2xhjslwxKOkevJapydiCOMdpink6gIf291qX0+99ai7g+VqUmYjIvn
7JyU3LAs5psubSJN52P/+kvJQSW/7t9iXiDLgdXyIYmakidhQ/fmqpyvre+/qRJycLBId4mi3HfW
NVjsWMmSkq1AennZDlNYfOIbnBoB9pSX5a4bURz1mozVNM+1SRadwHoVuo7R9wv5fZJ8zt91ahwh
PHW12iaF89WPi1LxUCd1pvNRnRnrYkX5Vxd6/EnMGxo7YvFo2qoGlDYc1rbekeO9wJHauaWaHmdZ
lx2JIKH8B8WMnD6ZNsk8Eoam0QV3KSVaKzkojkfBpShV0jGnL3qxk1AbuBkNE6d2RX4fquydpDdl
7ZdxePyiucEAvYnhv3ZEU5XAgbrJe/1ARowgUfoX84+atHZjEgIj6wF1GswRkK6RFxwWDWg7fmQ7
MNbkIwzGYuLxtE0qUWGCoGBybnU1z8uCnhGnk9Sp7GiHKxCtEs43YAeJbtqRXYNst5OGUtF5tEqg
XsXDcP+PNeux8HTD2sb8GmVCFes2Nu/8mfCqfjMPIGl0u9rEZu/f1wjJ09PI1olz7B6x2Ssx0b3I
4WKTPlYl25ui/SHH50M1471sGL0LBiICBO3m/fNbmf1MuyZNSdpFXYHTZIn7nqvnR88Gv+fxDfpD
Zg7R3UDVJCbALsVRrc2ccVfeU7134EQlCJFudhAvkAV9y2RPH1soVObjCK3BNVqZ+r6epQAi/3sh
OfD2F4hfILrCaB6TVV/pqWw783tzurzoYURatv8gwqlm96zKBxB7Y+MJZDUtDYuO82g6m0/7B4o+
mx45IOAyFHeMwdqbVwRF4oQB21Vw3y4vcSXdqCP7D4/8Qib1FYvxk1P2hVGdxMt//uZaMOoRhgQ+
goStG3xvle7yQJsk6gNGC0GA8VkyJWBlGI2QvqzRyUbDROoybP/HK+mxPiTcAl+jNiN6MtySB81Q
Ze9hdaWZOYxFeBhZ7+8iOJecv30/DXuJUYSmZ4ZolVZ/durePh3C6kinlPbuN8EE07ggvs5olmBh
UVF5CqyWKpkcfK0APrwA1gdP/9dOCU0mMxDM9Zot/DStLiB9n9JoNKPnBr7menSClTSJ2K0aGUWV
WAf12WpXg85yTMGc0fKoxky38Bu413Eq9BblLs/SE9xVYSiwVUrp4GVutzKPRNXEkX5+UbbQhWvc
o7HrC0sXjhmBMk69cgV6eKbRe3mZz36Q7Iz8wwiVrEsuF0VyOIKnVecfoe5n1/JrAViYHBjeVyWG
U4mMMsz21E93tXqwB/vDxD9xA6HkKM5ulMF1ig2Ls/xW4l1kay0XHouotYF57VYlmKCN0IlAia4J
ufhH8IkVBjFnpsWEPNBNDuHU8KfrRo3rjQ0ub/Pt30iLqeDdFZcQVpJxfQtpgTVnObithzq2ONuA
QaPmUYb/xnb4HrFs21yjPGGd3psgyaa10QiCcGquk1fEUl6nf71JW3GnPL2a7uI8am21OM+fY9vL
ZTGShLedikxEASAJTWUeDAjC9xbW7zPVlZMBNCL3fCsNBrCZ3cSAZF2Y0351lQpKaNZqkGdYIuCq
vgrSHIbefN0gUfh5VvTQYSmCqBOCyg6ChzYW/FO2KZ832xKM3XdIpXd+p7E48nhPHOaPUyV2M7MJ
Cnm1LRR9nkaxWSKHFlOtHWmTD9duieiQ3fAsm/c/37NVAh0R16wde98eFEAGKyeUg/mBZBE8e5sF
+riPb/Q5dkroqKFzZO7I2qHDj0j+bJu8E1PVNvUEPV4HnDPfprz97e1QPp8NFxNcJFfrFyDA5jzT
CjJR/SkH8O0kMrWpZNxRe2K6URPMTySrEIM4ZywbgcBviAIm+gyxsbraP0FcX0nnfvj4sjhkelVY
c6XL37cuCCbNZQCI9EmCfZOSCO0C4v301JAedYF4Pp7vaONuq53vWVZUgD9L3W3+LcjfECdtFXWv
2w9XJ7SHiiHDVHHR+gtLVImJXtwTgUbdrNPesX2p7dPbVPPHgZq4kJJ4b/Wa2cRF90FBOTNK1vPl
yc6oV5C5LUkHtgLw8quscEKTEVL81jaDjttmlzLmlKKL9OPvMazD6B586rm13x5W/BgtFQi0nxhc
31OdcTw+5M/MSbEFsNvTfSB3pGc6ZyDUNANCaVWCc/g9ErGlhF/3Uk2T7AeA0RaiKw6yah4sV/yA
HnaKNvUwvJJ/nCZGVyFNi1hcwGi/nKyrw8s65u3KlTZcooodzO12x0b0RZeN5NcxfJ4Gov8LcT5M
aGuzZM+FwtfQfbFvM/dhnqDvQEcLw8RZyi9JOOQvp9oQrPDsXhBwJOk0gZ8YWCD7iTt2WuKcoQI7
IwMzCSjY+/JC/XomJbWJOI85nIaaESI9mCjRhS/nUCMoVo6se9xtFh4dCWw9U15xS5Jj3TtQ/ztc
gA3gDLg143a/9Rx5BxzoWVXByq9wcu1bnY/Qs5O9t4tWzWIO5pQmmlet8VShfRltAFs+gtsJ67fU
RCpAAkvwaBAY12psIFzN0fvkHvUNdu5bAtnX92FiNhw8PGbpQVPopWTE8Ii/xEGk4wKo6FNU7E7p
HRWRINAVukNUyM9FEpd4IJNUBb6hXhZhrhueg7xOiGoHe1LsCgfWalrk/25VlKabJp9Gy9wA4JOF
gP5oluAEIlPSN+J1zvs9aiobEVC9TMtFUnD4JinfU2X2W93+M5fmQMW3EUIfvHdZ/3fiP4p1C0BY
ptLafAig2FeBjxw3ZpAzWLElppDiKHNN+iN3E16HveBpmlle6D7VFwniZV3uqHYTUxufVwJMlW+R
QC4AUXBTK6HGmynh3ek/A7myXXjOnTAIbY2UeE2yE1Ues0KlbLt7ccSlqXSZpQQyTW8WgkNLuT30
dWffFgbMukIRoyVJd4JMGjCNmNNmEKv3Wi4Y4jxYYUdwZn/EreoYv/9Z+eZucnBWd/fCbCeG8Rp5
LSXg8+YZgdsMDnttGXMc/HIKmKiYALiL5KyB5X7CSR+gJLEJgWcmZfQffL3m/kANpul7jG1+BeAi
upXSk8VmvIj1Kc/s0xFA4VyYKsywwJMck3wYdO6V4eHYm9yr8ZXZ83POy5zzQcavjVrwbuA4q2E7
5brV1xs2FN6zXS6L3FljYZpm4pa0cild9+mFdaOX/hQpVdBteZ9D0r9Dlttdd4zJuu7V4+u0vOmc
rBoW05YJ/Lhvng8Qgm1kBhHvuEqTn2yQPlo4IyYzoygtsgxntpEcJOl31DQKT3R2opkuWn4rwPWQ
MXDuB4jUImaZ8RPoyGkzT0pKgocHg0dFnyLknb+mrt+PNI+MWCPjfxa5pNFMJiaTcIehTfB6U7ei
3osNzoYYW5W9rCSTq6wd/CwTTBVU14cGD98iA/eNFJvpCvYmMKabGFYRCBHjVpHOw+yjTuReVYJK
X/Xz6r8p/DksDvVCN/Ji+zbtZXIwwZecJRcUBJoQAdoUR7Wo9ZwynBEvuxJfIWQeyRCfyVce5tLq
+KDvXi2TV33oGokS/KIIeHB71xQHiG8Xq5HKJhKj+qGvYI2SZ8EV208BYCU9YZU2CldPCxnykdUh
twwLs8EzhjN3dl2YT6Tdk/Tael3WBrz3Y5oI0h8nA34FSed09Dt16Mm85FJ+Ui/1Q/XX2qYu5jmZ
aftFR6Y8nCWS5aLAiqXMldqE/sQBbD9SdXmf+T6ZTfy2h+mMT3q8uaDhDEqEuxp3zgXjyshWzoG2
EnKi6LAtZ/hKm+zxjtQCrXx2mzzZIL7OHmISGJLTZ/5UQdAZSTu8rl8TKuoYbPtdPpZZQQDqp2Bk
txcI2n4+JcZ0t5f1cI3RPdUzHOt87UrtbhcXOfFjhEvsZQnopcRrtoyr4kiBCT6C/iJHiT6BM+GK
vnGEcbTlYZ4Ps0cb9xsbUn1VbvzlAMhm4ULb+rM3tyXfQwDYsauLBm5cU9usxBordTdcb2oc9At3
K4or07ySNiwW/tMVzvpid6w4H6JS4BJPSi9+R0/6rY964MN1TLqcN+OPagMPFMUDAireBaATxzPs
hjHG6mQdbAwaDHpsjmXJWINCXYcF4i7fKOwXl/QC3K1FQNk/MPCiKP1o+ewTO3MZ/4LR87hHsmNY
TzK++pEOrBjriIDii2/4EOXfYvisHoqKBBYtgZQRY67ZXKBpCqJ5xYYtzH8L/+Jd
`pragma protect end_protected
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="default"
`pragma protect author_info="default"
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
xI5rRsZ8D/mWscsXgMgqvONi1IR+WUmvlhOeHpoqbkmGbmmCKddy2Qan/TbchxUow2f4O04cfAEu
JYQ5L/DafoWEAHShGyHztGxj4EyJX7x8yqtcAWwgcJlMfy/2Z+sYHVx4ASnUNZeQ8HXpWibYIZuP
FjkTNuAr1SrdQnqwhH5cviaA/5OheQSigRQCP8RRQlRyBxc+biSsCZMpGISZFX2CZjSyU+7V2yWW
ay7r6zDWmMmDZjudTCI4MmCNXIWpp/bhBBuYrBSF+L/5EsYX/jb3bbE7tKSBxKDVS/NsrCqqNgPq
LE6lSb2eW+8BDcfgsBxnkhOXEUv0U/y1UADlGQ==

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="GoWin"
`pragma protect key_keyname="GoWin2016"
`pragma protect key_method="rsa"
`pragma protect key_block
kt+7rNkOSYrcXqbgq36Tjy1mVNbqyEaJJcQomY0hj5jTsV2loT+ykCqTokaSF04RFimKeTBrbOMs
fGmY0J0Y3FLdb9mRm02LfOxlSlD1IAUzPqmK1XSR8d/4MtempkKY0sPLjad2NV3YwFQOuIgbOEwQ
WJexgoWi794m/yDoUFziRVt8L8gAHObe8TsXdCCkIFw1w5BV4qiVphOfsBcAFfGjk1h0eqKL4hHd
+knMywKT44w7gE4DaneMKpcCfQ4X0hNR6jP67PdO/EqqXFjgnAn0wypmmiFT+lBYDb/eP0n/hSzE
W8aox1YjaQtyA9zwXG2XZMpfhHFKcSJlD/u2/Q==

`pragma protect data_keyowner="default-ip-vendor"
`pragma protect data_keyname="default-ip-key"
`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=146912)
`pragma protect data_block
RvX6YNnGq/QfZrX3+SpkwDzMRMPNyB83XtyOs+h+gSiynn1XhUeSuYChhjzO2tVQ1rH3F/vCPrla
hD6VUALEq2aW2Hihsr3uXIRTQj5xzzIbRGHkiW9zzagBUBHQ1t2CM3dtK6nASABOcV8Y7w4ecUgo
+FGcU4XD1XnCPgMKE/l6mkFBYJK3p4G5oqT6w/fkBvDg3xLScKDVq/Tv4x0ko2EZegEsdg7n2W6h
KdYcqV8Wmyhx/APgl+/v4ky60xtvtvxOdhzG9g6O/2c9eRbGVagU8j/JzWF/KZhoCpeaKoL77hTw
4YkPqcchCWCf5TJWEOIYrgLKQNHZeBx0HVVBONsWG+tPm0xV8jPkvAtArG1QvRgpq5Ou6zHO1uRg
x1W38QJXJnIOwo6+YU6f7L1DWvSCjO4RVHNWruN24eJS4RIr+GoHh2q4R7xeGe1036gtjRyFlG8v
CGj1DflgXLRxiwqsJLbkqIzYDYAokw/1aPxq1C3TGSsUHqAHdmFL4HzfcjGdHP55+kmCZLgWSN7X
UdXp0rg5ZLDKEMAeXNsm4wlX+ZacZ8KuvAIEEMG2Sb+ypjFeBQIteN4w0nDhQWqF8MZi6NEY49kS
Ip2tE9W6iGXAmeYPMNfxdwGDmj9lCRntPGcQuXFZsfLkY+07MWC83U0PUhVh2pxXJzA/6l5dmL/O
DhUtrfviWvu/kr4nw4Pzc/KCX9A5SyQ742+n8toFbgD1DYyQkc+lEnFcLx/FNuTS+Qvb7AgHmKBZ
pO+F/swanj3bjVISiu22AWWi8DiYVP1INVm5pzCRNe8ArJmhjb9HvTWOQQKVvJ0W5mfcTU64rgKf
uiZ65/qwhPpqR17Vly+k9OHvDTXZEhzk47ImGvd+d6oqrH0Wd8ILekrTMj4Gop/QsG68Xv0WfqA3
tWxpJ3bwym7lz4G9QPRHsP90e79NEHGNSJgwOg27yT4N9m/2qZpPqEH10o0bNDAOoY0w+oFFsHeo
iK81xEiuX6aPLXJ+1rtOq8d4gDvlmAxYHovvVEHXouDFcffo1He8BOoMcCevG7mWatagvywydgaT
kM3pNsp3r+qVQbuRMxWjLzeXOCoaDxoLjH2uTJOVCjSSxTf/dcmTWVJkwnnW71J66IGfE7UqSF6s
aB6QKiVLsT2q4nsKFX9x81P6oSOqwQbi0+GUWzt6mIyOArk5WG0QoJsuLZvJwbjVYzGX5VZSHG8H
+NgJtnYxZY2pG72l5qJpZyYtwV7b8QIOwQu1Y2w9+GgUlbr6iTZe1FheSjLDJaByxz6VJLYwQjMd
6TE3wHJqeCXKxALmX/WcoN90l56TSE/VCzSegUVlX/4dszbW+HnkYhlQlugdn2LyC+Ls7FpP8e41
CDL5xw0VidoXMFICj0qwuXUqtgTr4xpS2DfsC3qfS8aZWxAK8x4PPKHj8O5d5wfniHP/awR++5k4
wUEHoCQcS/K66vtPUWq7Z8/OG3VW9LGKYzEykYB34b74AD5iTNQU9ee1b/UMg+7nU8ZNntdvC2IP
G/cTFgGgSwKOfjJfB9lJtgiozPxCcKV+NlBsYt9f+ciL3TgpCClZ2c4oxxAlpImMo9MqrpBoRHAY
bJtLhvB42bX6yIIJx53QcVY2NbWBDdL5pb5INLfE8EtV7cBEB7eeB70QkwHRgXtW2m60aP1DMt4g
WBlLRzhmbTH3vxmzo4rjaZ/NZ2skIUNuSdzJKbWqT6gWSpYbFQNbwtxYqt/Nvszy3R4fSrY0oFLU
TdI/9naCEhfehhNAit3pZgZuglbAAVPmlbwHNtknDFkqhK0LFR7qX19ueCgNErQ95nhfFMHkwbax
kw0Jia0SHyj5AvoU23KmAXEVJUuUzLJxH1DPvLfl7r190glQPj+W0n3fl6XsbFeKhtbt1ivQNkCd
xoHrK2NqpXfuh/TDBcRvRMUYJiDzrgn51Pqpm7xvGVcUez3wJPL2X3unPl//3MARNNUAjKy6833s
qnbYlO9vxTC6sHsOERdCqtPc2vSs4edmS6Jg0YMRNN+RGIFJL8ANDykwDIvPQfZd5nKUZzyfmpv1
HlXPKIAUBO5Wcpax6k2EXjKqM2GY8BtQiJ7hIzN14vOQXYiSQ97pape8XdPAQrdpFwUZgWQp59u3
6uWtAU/UO+xPK0m0ZlPNGTSBDNqsgoulu8UgjyxKd6oRvSQMZ5hUbrBnEhEvsLb/VdVDKwfajbL0
OJW4dwdaBa3cmEhoHUUqy3P46WMM0PKQjhdrpsHkK/vLPmNRvcysY7GNCszogl4ReNeRgvyzNxqu
FQWVOb6IYz0cXFDz04aiuMXFfe00I7Lm65UAW6zMTLlbwnwHYCl+WTkbPcQluMQy0P9jsNb8XijH
xZBEDY/0XSXHbeRLeqAYIGvfaZ5tUM+0bpK8c+/RSRe1SO5k6ftKrnXtvsNGbbfS/3DssaveDJdk
Qtq9/CLPcRpipOs5gfmmcLr25pol6h7zXrxGOSFWiZW/NrL9+cs271zojbmYBPXuGa0fWLjBbE1V
l3RC0IcLjG5YfUGWDh1BHb/5OGGUgkqYnZZanBJNw5brT0F3waxJba+yt3LuNTHOLAB37XeolC8f
N2/fJh01bYoLcNKhJYet/3ZiQJzw2BkDvIDSOMKf+m+5gxwhkduk7W8IURvuiycVeEjvT7Y4B35B
Q+wx2eHeQZj8I6L6RU5z5sTiboiswQm343r3Hlv9nJHV3ndkDgXGAvNZOxQOPWjDd8Iq5jd3QFex
p2kbyfp6KuWV/ZMKB9iTcLXMUJS0fHuWkUHnz5H80TXPlkhFoFGdGXnokmtKxj/KcZox6ef5q4WC
H/RKJKoiWx0Qx+uEor0jsdVPjJNqIf6o8/oDjvSXgOzz6B1EP/gzP6Sxo1N1jDopIHb9SET77s64
cAV1U7yC8uq4r1ebw+OXgps6W9PiMZjqtu8jIghj7nwzclj4p28vtIcHE5OYBfp5Cf4EIg4veOCP
gYq2wQhM+ww+Y1NkND9tgOJYYdoj+ZWLzjpjHLyEwddfIRq0yiBZVN8bnfZbwMTOQcJcSej2oAE0
zSVceOWfzN/7u3Ysp6kEYByJpj8VMpWqMF1tuXMhYBw0+Lpy9V03uHJV/bKpa0uoD80zEkxNxKhe
cvDN0NceqiiJlBKfokvOgYf4oE1E4TCttb0ype3J0RHH+WCEHvOOzURd7qldx2GC3iKNRD5YLWzK
CQ3teBLkhSzNAausskhXMmxNRy8Mh4ihy6P4EZ6KsisLZCp0wyezRak9MdNbxVviGHTK/ulvfH34
63fel6CS6rv1AmQjxeeQm+OKESbJ3HiGySyvQaMhDZabdjqiXj0jxSnrbh1YwrWmD2zOM+W9Dbmv
TlnVk8sKJNl6vv4PloRIbETzkNwqLin+WWty2O3oUrhPiE9o2slVzqQMPE64G/2ezd0N1VoST4kS
C+Jf0ph7TZkmX9DECM351ULYXjuNOp4Srp26776fLRGgCEojCZL9EET7JWsDISTAJEam+S4658Uc
kz9Th2e1vjPTM1vPEPF9IOfvXoX0rlT+17tOejGAUA9iQk/EmfhTg7u0SkOHQzuCDVJgSfQ1hbmF
qC8eNQ/hLYjvDJm2ISG1gP4LgqZ3Amb19firTJyxiMm8axWP2HTjxQTllptqxfIJon1luSRjp8nm
ESvd2jGoWgD6GK1bgJMBZIar5UqjxvDMDzdsX6gQ7Nztg2DwPsztOd0UyTPvjsVzuZzr2Kd8ZdIF
tEUpe6W4nJdMFRoTKUMSFyxcpvs1DPiHiEhfplEYvy+MkeJ11Wn53MchOreQM9idnBXnm68OYv1I
ndImGAxHCwYmBAaP5JY/ykKWs1N0UX76IBiYrNgww1Ww90vrJKd3K9ArbM0HXXYSuw/yzKNNxoxw
X4PaqGaF6WYQT3bQ/NAHMWThIQ2R9wG79/pqagscepTu3nnuq5uOZRTyHJ8jGU79NQz8CgSi29yh
mWsS46ASu3j7MPLuwqHd7bPnJ3Bhyszw56XJwXgRDI/lMtZJph7UzeAw7qQxmzVNdfutW7Gd2Pny
kJa7pMAedMTkbheEcFVD5NSz1qO3Rg5XET2Xm/ngrqUtaabND+QusnXDdFBSgejWG97f12IVF+LY
+NUwk7moq+SKdJvqMXPpCZsIHBusMrRYPJB1zZNxPEW3SZfJULk7wIsEWjmqRRNFzBDs2o5VkQI5
5WEtRm4Cthz849+G8TJOKfgIaRugkRqUY/0lUAnGbjyyIreQhT4A8mQTGpYXW2W+YtA1z6ZdbkNZ
kpORs2Q1PTiuhRTwUOLf7H3Nm23HUJgkr20jhltqJX2UbdJMvQMo9UiSX4n4MsCSglfzhg5XljXl
X8AGZNY56CXxzijDIDMC37SoYa7J5WfIDzGq5Dj/tIealDHMGCi07uCqxfz3GXqvjvKAFif5uQDt
vipgsCuONqRWzUU0U6tJ+3GgzTUzkwdPQB4zURHqoA8sNMDaO7HWr4rR/XeK6va+2IsQgYPgAS2k
kr22YMag7b3bn7jSkLzO7/iBr+2fhdUIpZGRInbG4i0lnYgqMGU5XUvgwJLGWRxKdaPwHanqZdyB
Jtui+sswx+OJS6IECpwEwU2p0h4QqJs7wMAytle3DyS4haPI+Ib1HdFasNHILBSBySFfrB5tOYVy
yjipE/gybKaquAjeoBb7nDscmY6tfVRH3EkBFLaVrhhMTAPcKJyC4vxc5zMaj9URcJlREzLM6a8j
6zVGv88TWxh/HEPduenhDuQn5Kk+EHblSN3pxH9M1EyH80o4XY0W5HoEpvN17+nqavwP2oRylHqT
Bb1IsKUpYt2lUbmWq5AQvCkbMqpobZrlsv69E5b5F0OniUyUYv3BZ1a9yuGnRzIthl/0oVkKMzcR
irE9w5taAJeHHIR6mN2YE2q+I8LVpOEn+DUtef5fNa7DIqIth/Ccr02PHooKFLK7u2p7/BaH4Tu5
M4lyaATteRxmSgh8Y8b88eQB2iD12vQ6+2zDGRX/phZN6vCjcMRtnZJ5MSgXZhyLPOvXjNcUIXPo
XFhOSaZGUjCGVIDL55bbJ6nvl275dQmb+iq8QTSBoVplXk6p/CrtJ6NoQrDUx2ayrggcLYXnjJ+t
caImRX5jEhymqBLTtgXQ6iMlTiuH7CeoXmuNuE12CDDfElvAvrHsugf1xbZMqJA8s4ahsTSFBgF2
8csRNxJ+elG9GI4F63K5NsNf20IwZlnkkWkRCcZ2HrhemUlVBieUgLDKM8f351Y9jlEB2g8kFSat
ed23HeSvQnJR4JoY9VgSr5tH88zg2pJsaDY/N+JAAiPKpt+/irLEtO90PzpBC9R35OjzhF4CRGyk
PUYpnyYu/hRxFBmwrTAQUKucZ2Bi5ZYNXWJ+t3ESXB/OIrHLF2gxU/fSBf5OQaLr6LkLafSEUFNA
rHBD9RqCUHUavmtZDuQcF/hE+d2gM4r3Uly4X03rZr4+1bpGu4dhKvxinmMqPzovPQ6AF/H9jNT7
5L5qZRr7xAEmRneyQutdEx0bUUuOZhQ/iAvM1isqVsyjwyKcQ1ZQZ2Ko5FEmZHr37SBwEGBTAH9R
dm1JEv/c2fESzk79Ca8j9eSDcEifvws3wL1El/LEZq759oCuaFdkV6hAmcn+ATc2ME1WEZwo7VTk
KcYGHJxxRtofJFw4s5rnBwQs4aqiz4GhhVEuGjfaoqHG5smaTRHDziTc3wtOppYoO9R59jbse0c+
7YuJkGpNodRTrUevAfaIPDSvebQoi+77Wr3vJ6eOVZ9pCnVCY5SMFLGpGpZY4lgdfXyrvRvir7Jx
e9zCokrxDtBX+ZkKktZNO+J9flqTJkNV3GreIEcoLtOJ5V+DJBt4nOGWfKAxuVDqc8sAJZmeSLUB
lNeAKtA9Q41WU5tJNRtNKIJjXxg1oVat4XaQkKP0UrzZQ9OWJ/UMrd9r04hr2+C4ZUHLrLI6KBXM
XYuWSe6I6nnpPc27tJeSi3GhYNaUZhAeZUgFjHiAPqZZR4nmHQmljzezyxqCnXlO/ioC24RlNWc9
67JUgoMSEmRXM6KUN/FgCqsZZNXpOBSVA5LSwUwPi0eGYUYZidyHwsV6WBGTLdH9pwG5USVOU4ZT
XXWAfgnv0IfF5LmXSgG4anyB4oOYo38sELbHPfVMRHE88g8hQ6Qfe60r2Nq7fqJ7bjE6SECvdMxu
vNY3fiLboPg93Ewgwguvu+dOoYqQ4XeqMJmcfCKun4kG4E3MMBd6E6aPCIWVKbMD4oCnsJLwV+ig
wYlUUWDXWbHJo5VPAcPTDP6ErbG32uj71z/vjrvTrurGIwZMQhhyiPyuzA95uPxnqJgBnbbLibmc
SZVT7BWlwni3Tses/d1swXZVM6g0dPq7P5iZA/uRAlKxf09plvCQXlFzn8t/cuj+k+M9/bNa9gmx
/jBlYZfTT1spoJLSKpBAWA8/FGSVWbNYi5q0JA3pB5rUs2WS1DOd+7Rkl7p9zHSQil0Y7At8DCT9
W9ZBl8fcl3btxt2/Nbv5c6I7+UaPtnAnq2PKRYDZut6IXC5U52J3FeNdhGwc1Xpj4tZb0/Qn3++y
nRp6OutdVI3pEZL/ZvkP9JrWex8mraazcaEvwzN+T+JR3IpaAXEWsJUM+74LdboGBIxpW5XOA8NO
aqS5MzEp+SJb2iFuGYFac/plG3ZhmgZmWn97HcdS1CvXYWRJ/svXAdUOSR92+HkpNsJbNOdgOuqn
Si2Y12z01McozfjCWbvUa6u2ti/HmjCf7BzAQHyp/MY0dXUb9R+qtulgBP4+w9CXPYBDOSn6pk9R
0RSU3FyrcmVTCGlyVqfd+FzrR8B8ZuHddQ1NLL0vlMb88fr+D06v7z2ZIdQQqZkZLD5Hl2kM6LkO
WwZds9Uf4RR5YO8ZwL0EF6mCNR/8PSdlo0DYn5arIYcLoEWsgKD7mSpaehJ/8JPTV9kxoJg1d49e
FpGDznkkQ4Na5b2goC/hd67lzCtG+ZydH8g3O0uSV0Us2yFsMVYjg+3l/aZ43e/sPxfFT0ykNpU2
lkKhrZxxjzsCtk7ml40+hjsFKtU/kgvj2ONqDXlOHCv4iQ9NdZFtLddyLIFUl0Wu7MfWSljgTjJ3
wQJP4NKhsNf3Jl9qcL0MDNaW7Bpc+/cI35AaQjsjpD2CfB8ojqkFTXAlzQYNG3i0tcke3qAmdtGU
CSoZcxB3g1MuwPlnq2eFY0warhJ7K09DiIrtO8sSnKW8yhR23PfBRFj4qZTt5LlO2v5gqxZoovPR
rwM7Bcf/TxEO8VlwIs1xXDTB+0afVWClWHUv5WEOC5CmUY1tk5qNtyPw0M2CVU/OxrPyvj7AYeD8
Cc+QMe+wRx9S2Z67qVFHIUjHXDnEO50gNHxxb/YNTqEQcjP06NN43jtTNnheInt22m/XLvZbIY0N
5DB3VjepUHAecfHWpzdljmnCZI6NkubKv7uVGYa01ULOsNaZt0p8lbrwfJsGQqLdh7wi8GUTYIpe
pEk2d8rsipTWrkWosE6ZWQVwD8sz6k3vCm6/uH3UwcAiUBDNCJh2DIAI/z+SXDKCRmCP4Uy7xct9
XBKukMW7X1krNcDoaxaSG04GiDQOpa0n7di4k2SXryqD4Cu/T9MecI70M35F/hTk40/quE4m6Ilb
s9+umDk5Gs2TK2cKTUp0/+rIy6L8Wzqo8RNq37YDWl8JeMFF6bKSbFYFM6G7L/gk7ZIeFhoSYNMR
LIgkp2iGhRypR9vurkTG7eEmiVB/WKkj3Ig3NSA2JR8Z5JHnfAVj5Dghs8dUvbPus8XEIhxcdJ0q
3LuD42IdkkfsiQj5+H5eyEFIWNfHgukTQluSc33BtfugeWSJc8sn1rBRG2HhNI/dBPLcoeAl96qT
pu0rITg4msI3S/IQ2MkWYX9lS/Ta0UdUNgGjE700JqWAiK9ZY94mYT0XNF/6TMbyEgnAiG4PxjW7
2Z5rkBGxH/HfJICTuykO6d7d4S5GmoMfCZhjgWb7w7dc77TxWDQwj+bKuDAf6SRURheQnFOTl5QC
DyoCwqaK4M5S9CzO1Fs20ZN9ClrwsLJtT1Z89WNsOgADtMuPoSNsCStOj2zY6041ficeBYGi4bm7
eIulbtkjyTvd/mxdGdP6UrcVhFGT8Wx15FSKSc2mPRBROokvmqhfMM75tFYM4AdnfMc2UrYRaE7u
jIWKVa+44FcTjlqOow7nwK0ZedQg/Ss4eouB4MH3JIsrwDkuGEKl1hAjCsfpBQlPKEfOjmPn7mf+
Q/jBcz3N0pCaPAvGahN7TvEcrZc4YaVPimp+kg7vXX4RHhwRb3nQAU20c/PTTdj5wAn3Ur/pO++n
NJyk7Mle7QuRPZV6mrRvuWtoFWgrMgVzGxaU4hzkVwxDTY0Jwj6SZRpTX+Ed6P9RfZZ3Jh+nC8Xx
g5/6SfRJ/230rhiXDobDGSFREq4rCyivGPqEfrIxlHtakEeWWW5+hTvVEeaoX8t4iJVPzMWSLNkq
mw8mhWAsUXLIxRj3/s7FkLW4yHg6ET54GaMyEdiXFgvGT2RO95+PUyRlhG4QMo/TZ1T/OAcbJSBC
GeMGV/nwF4C4k3qi5hkR2JvZaKfDdCEG9WWx+eH8O2uaXjdQIIS86pn1HmKdpjLytblWVhC8lD66
mgY2qXpQbaFwrIgvIWZhfeNf+7iZAaH+w5iVLAGcuBIGgNkzJcEiULqbPP/xLWT3hZwn1rXVD6Nf
VMGCnYYa/y8N5THKHAgj5ob4ugLsxMQ/1nb4bD4f1NclLNuGYAfDFxV7Bbb4OV098EuisOWy4TyD
pH5/25njRbPIjjzEPYFw7UmUik7vim30ycNtjCvprELESleTNqPkksvFyNWRrYpeJBLNAA/pblK0
BUskMF5bYVZHG2pHApn1uFT6NqSmAm/4peYpDDNa/1s8kl961WgC/FW7LhHrhEAjt2QNBlRHo4nz
pb8quR6u8GU8VH2AM+AyVm1AXB3KupszzysJI+igbDkjE7j5w500LH0xFrpKy8MzRSbGimAg88M3
bR8zntZVVwgCCUzjO4RIUepJ1CRlTtrtb1Bl6Lh6uCHdaCbiNQvWrxOBKlgApx8PeRbfH4jiO9IL
hp/6ufNwT9aYLEHRkX+4dyQLZFAnXVQNwlZr++Jc7eSUrzDCH2f/GG9LDVQeZo17EvRMUy8ysQam
RJdKFnPQXb2GQ2YjuVR8DfPhP+b0AcJZIBS3bfjN+aOsiP3alVupbfr64F1NnY+eVgD9pkV9Fuc7
+AOSCrkX7hzt0Pq5zN+7DPWNqBHOZufn87yDBaxGgnwlQ+ptwLfGqvnFPZWpL5KOSHCSqiDMtJsF
4GyWm/BYDd4aSCx4wsEwHT3myAj7CRZHdejRiQXpol90EdGOH2QbRsf8/r2WY2wT2TNQYOmPOWwj
NxkTB4h4P1MtutTFmFj8VPT+lE3HQPzxg7fzNmVBYH022nuJDvoowLZQmlwuUfcBhS/G874xIrA7
f2DO4q8H7yZVEO/zgVWK0J5sd8hWCdKdCsiOWiWue2PvLBsw8U3axgItKU0+DLDhqA8Jg3rrrulo
yYU7BAyTZrt0bj6kyscTXxD2a7wjSyX7xOkE3aMATFMlsmOGGceH/ErXS+KeK/t+zGZl3R32ByHU
tfMZaFgWpbgvmgMLbO59zC3Z6kfXm9dHqB9ayYDGq+wQvDmb6WKQsegP4XnfmzdHjCU6q/R0DqwA
/bBNSL41nlEC7lDsPR9S1XV1DWAZkwWFITIQZaYlhoXsiroegFkOkzAaOLPyef9MQ5d0NwZ9dOst
LPG05IVNXtN/oUU2IYl/652Ycivr3rXPt12MbahsBReOQ4QLhKnZZdlEpm8UXqAi91lydCoB9qV4
zJnXh3729W1GwN0rT05d2XJKaL1AEG09g6Qd4SFjkCbp42qdbxPZ30G8rnmRtBxzmbWu5dU2Bp4/
JjCJmhMMPOI9K2RQ0CfJVJR04eUIhihhA9ZObFJWUcq+YSEzmdjpyd5ULb4JjB5Xfk0mZ1Feo0uR
6W3l2G/Kp5yNcE6BeUqIWkJUC4CHEikbsfVSMvhqmrZRgr3jecjTi7BI5nhi0qsC1yj6WfvRyPLI
Gb+/PCLG8JeFbkeo/KexqKscv3qsHNSG0im5ElGYZsoexn4i/WsWhUGG1BUjGg4tjHzJTe9cQaDd
vIEk49JcMRpyypo6iGb3sEiSE8heoGZoYSHMcvoIHheAi5O8gqLFrHALbJcIZwJHmKpdl8EfJQDS
BgBrsKQEWf98cjNJ0SnsQg6Ol9+CugVGiytVwREy6zBB19b50OVc3Rsfy6eJtAGYwjHsOg6i0lsx
8ipvdFD9a7o/CXhwxRMfaXfAVN0IQvGQe7hlPjWIcX9SsVrgM2SWXGlVJbEkNfXr1S789AxuJ5zQ
J26/iptYdNksXHGD88C7k8JZwycy2MpnIdoFiH0ifWQrBqLKg6zo9eU/40Yke6iklHK8KlurF5N4
6Pitlq+G2t6JVfenurqrlwA93LSV6ox5128glGOX0SDsuK1H1aV0sjn4O4NihN7NRUsuKqOuINky
WpMAkfXP5h3waEnQBrwDWdDY/bnK2JYNCQJmmT+KQ5zvhNYZ2ZfsNXAhT5XU0C1Zgvl/Uyf13cgP
c6lwwxniD/XbpkD0soP9Ya5yaSYxEj5kmg+jhP8pw5uswRCnSwqkV3BxO3M6QjjH8SgxDa+FU5Fw
QC39uI/+irq1qSC3p7Tqf7tTGnmG+FCV8zIIxILgrC6rUrnaONjRc0MkX5vPg94f5gfuBazqnB1s
Qg+wE7CtqHnsGiArFXLk6iuQdsoCcItnTxi85SKQ76ksFkvsxYApnrHCe3vl4jc+641S/ukxqq3Y
GeaQ6A13eWOeoveTZgJzhLyCB4c3ObMvBcvSEqGK434Rp7P66v10s3Jcp391x1fZ9SD3xvfYzNr9
OgCEbMigZiH2dcEDV7zIOGLzRbwiGLRPDCu/Kl+AnTX8dFwl/eNrH9GUyq2SEaAXEUHnv09BpbGJ
EKyChbzTNOh3CTlTbSqpAGmpVZBamMqFewlotxFf2jEcNRqNC3PhYYE5p6mNj8pH1KYZxlvxPZw6
AKcQ0zZzJwSOg5jDwrWCE1DiWkHmS3r5JeKDIlTE6sJYSjqTagAnSEQK8wcJbpeyAbIEu+hd7DoW
1oIzHzO1ZxAJUCLt4ApncTWTUkVuOIBWIrwCwmgaXEQStyLMtVvdmIW9lOUCbIjwD3KlqVTDHuH7
0U6Nhbs3LfVXknC5Ge6NzuPbggEFBwbSk/x0qwV5tPD3RsFEg6rQ6yV9sSuYEacx1mRDpMpVeYLq
h1/0Td/UgLkz9dKI4SqRLxG3lW8HhPYLSm/6uC8wZ6gtfIAXzZ38mFNwDDzHIyhgd2rz7K9CWOZn
242152v2870W99aCl8641slMsHeby/33F6NH+3WlXyd1Y1eC6iRLe78SwOLKvf2MbTK6Xe0JwIrH
YFc2p8dJD4WgyqTIgOIEZYo7kUpi5kqyo5zyVWBFLHGuN6AGgHdO8P4KPMhktUfTN6upDdpO5D3u
LlXJJTBftJmrbsgx7peQn1KFuve21niHbeqm0NIK/t+ceYcS4PE9RXTYO72RSTcSUqwtBTHoPq3S
jTMnM/5xtbN7QWcpa7hCdDZOTANHWEJ4FAapmHgeyHJZPj5ut9ZO+OiL2x//O18DZSqblhPwQ0AG
LhISfvMe+eH1yLtywX2MRvCtnek2h0wf1uC0rgXPDytw6lOZ2LW723VMDgrhHAVfWniqo6u6zSW7
P8YdYg2agfm3aiNoGgoVsCBp9AQp83hE6CN2/Tuld4t9ajXQwEo3zsTijGqdUlD0rBDNn5dfH2YN
Emk1FW13RvswOoHq8JLef54my3oH4cAvkenfsDJB+J0LjKxt7l9S14TdIevC1BYJIYl7Lwnyt0Ji
uVF0niYXPQY5rSIMdXODnZzKG6GJVML0+ur/nFbEOKYxvxoDgmOmMdRVdfqNbRziI6xs+iUOrBut
WGiFaTMDzcaOmaEMxy+hMNJIaMytvYqVeDRBuuZuv5TwD12xdP3bsr5PA875cU/wmMw0F6WoPuNY
/BkZwiMfVKWjd6lb3BKuqyHcb3OpDmhNcO/U1C8ivmOCCQEK52sZEVQYSKiw7czNeb/hfB7Aqug9
v0gMcb3hqlkSfTr6osmbyy1XWNS1/jbPw30X3cpgAIbdo48NeogfDfN+0pYUUyINKS51hoehxD0v
wxshDVvrwks4aNJcavIfbfUj8hv37J99quOF2bOCLkIrd9wY6KgT+A+pkon0MY2nzUUj2OCecw4B
jPGpIPLGhaLeE1I1mBzxn2RqGdycHod5/Z/Dh7UmRuMUEO7MStuFg003rByhXf4h9iHYYNK7pMux
e5ih8rh8jaiQbFP7kKMGK00bXCzZj2Vv1dUmrFVwokEIgKItkxGI0Bpbg3DIcu+7nYX6bA8sMTeg
v/aYlQYsKEJtpPUMXq5vmU4xEAgNgTAnM9A6PbFkMfM/wmvDfNq+CjJXJ/xcKcbJB+09vBKrw6x5
9Vfro2FtwgC93y4S8BEzsS2e+AjtoFQK2eo1EAu/hAvrh+F2suNa4vnDCkZ+vk/BLffFOrwMt+yg
5QD3RubZ8qxlFYsslh2/bSuJDPMkDHQSDxDg9IcIcqbt1pafMN8tJ8bDE4tSgAlUJchcU+xCVdgh
T6VUZ93fRHKNQLj5SB0fwgf7vTAxKuLod72LWkOVlQtojnvAMo5PirRrdSkTjIsvIy6DaXLcXqVB
ggT/13buQgJsmJC8uCo4oK6JtqDIQa35q8YzD4Eq/6k7NDUj/u2J7wl6kh21s2NypQ4iUBgteyE0
+M/QWUlFYrebPEpS92j7Vi+So9K7PbX9FwhgI2E74blwaD+gqAX+4q0QPk/xhB/K71XXZCXkT0fl
qeQsZQbqJ1npoPM9vDrXik0yHDk57Bu6+O1xy8E5Clg7sk7NWaMLiQCS8AsRJxzU+yRd9NXx9TCF
iuvFxzbhWcsPYsKCiS/wRaEq3fJ4IinHfTqKROEuef8GUu5KWs/qK8vmZJXWKRwBe2qLaDT2uw+K
/a5PR2Gd010hu7iefli8LSdUE0M4h+1MI3kb7F1ukuIENa1sX7rTCFdTPQMzEMnVxudVZHO6gglF
Wp2KuWlMCjCrX2rF8xeKHh03mQxH50BlM3np/OZFoDb+WGrkpT4o9GXdJkQGF0TZ8kY7jYP/Of4s
UPyiJli0lPndI5vN6a/q7IaFQspWHXjJ8WjKXpKXJJ4azHL622GCQ8AdatoJxZjXFpqYO/UF/dEC
2s34/hMH1TDHrfK1ML8QrV6Ml3zoRK8EDKUkpVLaxIC5r46szv+NxeEChr4ZT5CGjweEFC0o/Z6s
8vSH6kkLECpinYyC6oFSZiCSo/lhmMr/n/vVoXDRyCejed+ife2h6C2mbHiLRNiGUgbpqF+plWoB
KZu6pWvmjrz4pOHXdm9SE+wP+T7lMrsF4iIAQQ1IuhVfiTf39Cg9onWkXZs8xVd3sg4KCgGLZaGd
dIr+MjRtRy60/ceavgMbE1aUw4Y2Yvdgf2i+eb3gmQlFqVRipWNFSSQl2YWmPQXMwrwx9KUscXqi
dZqLvF7x4ULrh2eibblQYM6Jy6bdDjS5+YCk9VJ9MNSiOtrrkrAHWwvmN1OzRPsq48HXMgXcIWVZ
/mwrs0yp/u61GiA90141lMZVX4AgyCvbD2HS2ACm4DC16bl+vVbdi7W4X4M8PNI55E5Q6Jld8aB/
vXvd4f64cXW1HGzhZaqtNtcj7iLKK9u11WGYk9t2JwW/0fKmBMIXMLYNRQmMp/RJdxSR+6bbP5/6
gJY2g8j1igHSDYw/7aErc70ZVEHEm3hPzjqZzFCkTi+VKfuCNwcCN+UrvkdKapNQoVsDKHEv0VuV
zaCZz03yxpkDd6+1aPnDmndKzSziz3wWelXqyRf5jDkdKyvXGXFW4MDq7xA1W6gVBjkD5yisCY9Z
Rf8CgGH0fy8dbxcShfO5/ve0isB8v/D+2U2Gs79OUZCa6s8v2KGfvVxLLHXgnb2cunL6WPhPBeIK
9kcCpte0WysQVlvImcL/heXxCXoonW+Z/iXQ9umElcJVkQ9nNKellnZL9+GjUMnAcBLR2TdrwG25
RpHm8DjmHiqfQ5I15DUUKA/XxKLjhjYBwSlfrFFWYmwiGf4R0Ot7NsBA9krPt9+j7g1uPXi0OHTv
qLJZu/nh8cjQ7+9NnIikzVY0hffskxdJ9bBdd/0wVzR9vH4hlBuyz01N43mx4s+GA6Xo5iIOB6xK
m11XBxv5ymyxnk0zniFIiVWFMpIaL7oGur8HdambjACW7NnE6NcA8PhEjgPncL3BAEDMuV3t7ipB
xvyiBeeuMAY8bsAyibEAbiKLWHlid9Jv5sAZUYYzfK2ZkxW0dOsMNN4BEVCxWH8StX+fECtwuR01
bq7oJDfvfZ0dfT0EfayqsHtfSNLlH/Ab47qrL4D4sNTeGEiK16Qzdo124T4nd4VHaf/s1cdEppEv
m/aMF7GCP0Yz0M4VKdM1mv0O/R31yuvj0iwYfzpfK/mNkzTwzUTqmvLTbSmMxacbg0oDMhQCjBSe
7CCty9OT1kyBpLTop1RZAQAt2FKX4xuZl1aPmJqX14I+6GiTX7yTiOOUEWIXMTMCKjKMHX0ZZ4Wd
WU9JGw5X4E2NJ1/Zmi0t4p/oBbylhI7/a+8nIEolXXEiHy5oHRR1gH/JIjBP6n1QdMi1JEdjuQiu
XuxH0FLMw3te/9Da9wKL2Z7U6PpInCAkJs8BPBKEVmet5EG6eeGk4nPg+spVt1Wd8hqcX8hzJtP+
3rgiS8wHCil0nqJ6yhN/Vp38Spnc39VxasKdqRkXlsM9dBy++o6vltbVBmFEmtZBs/V2vEILe4L3
qTx8QoKgzFcOz5jJEVn7c56hUUGUl8mjP7GJh2nZMrMlX1iln9SbeAcrguAV1WG7tOadhBmzkYw4
wk52CWmYtR4fE+FGl7i5F8l9+EiKWo6rSWHVSvd969KOWgXTaftLKSKd4YytAgyhZ8LBYusFdmTS
MK+sXKMVmSGSZBUfeGDgIV1CVk91IPV0wIqXTUfrnR7JN7kSv7yHxpQyI1RJBrxFgvS83TX93BZI
aKfh4d8RCeNAyeeamqqHs/7UxwxAqvdpLJ5YTJuflrQ38wwoBqeWp2zr8f2TNvTTqyb5x3IL+4ir
6rG5sS0IQR5UlceWSSDZxFA3tpNKUsCCaRgYFA5lYwhsOq19ngw3rWMV+a3SXRJI8l9mQO6ZdGIz
O9q3C+Kmo6Jje7QMwXauJWrKXvq72XgUxJV6ih5nBJAvgAK8JHF00VCIsY9Pk8VQ+jWxpE3qwQ3a
taZqaHSJqqdsIol5lviJazUImps2LilAJBAl0ATVpOvI1FiyS5HDtbB3j0HvzBeNYBY1M1fG6yw4
aMzD8OCVxXbub+65jMbybjIvuUuxYp8pXnTiJoDvAyw+Xjm2yNguFOzElZGzYekaontAd/cXGBrT
5/Zw3T0rY4Q1yHyXDnX9+OXYS/SoDq3clhTYEzD0phWbJRxv9WkRe8RRAmFHi6mN8yUTQsithPp6
xwtKb3SXTaDtw4wf8ylaA/F4/o9h2EVlAlFn27K+oElBI0VhlVUodqyBIIW8UGKZ12+tYx/0z54D
pLMy6At5s9CxzeTH2BFiHkBdf/THlxo/TzeQsCEMc7ZhfBDAdaclK7mtlGKEbBY3pytQ0soW20ML
mfrFTz3RmH/42HD1/LAFcaqmYzCyalLODAEj4XbP+M1ws7papbS2+t8fnqYT8eooJUEhgpb1Au2V
x2piPxYH+PXBpVvPfZiDNDUF2c8HPfFcGcEZrQRttaBRXgAfyjkw6FWy7ebaw4Q0X/xKBuJabwRO
Xc1CdfOPBmkFXhAcNyAtUatYvfUYS8E8hxnXTCC2R1WEi/7rermKsfWir4cdjwhnYNPnCYEPoONd
g4ebT8kc73YYPj8ylV2QfXkrUfOTFTORnzjpk7AeJ5E8GfNh/Yz0X8DVr2PYNEisdiQIthDY20ul
2EwPEiPDp8IYcgkWXbBbT1WF9H/EFpa2eNdUY3jwFRUFhNbKljvgwB2rOQArd6JLr/emOvW9aB6t
cVuvEmVcf9tyGlWVUixamwxpkBAIIr4LnKP9G8ukqKdtn4tijDD7CufeEhA+mA7ceTjWdZwysuSI
/7DaGXwDiE13q+uEQU2nsLZfGuhVTm7kzskWiwL/KSuHEyZrh9IRkLBaE0tl6eWH3QzuWAJmvWou
dHiF1VC6mqE3NlnlEFYIOWIST3ruYZP4DweK4+2brmRn9C06FtGAQ2G9e4QPa6ZDIRjSMHSBVmnP
wkqXvMceD7f34/MqzCuT2XhtlRDOpNgUSfi8CL7TpgnHtYpWi1/6XzYkAJmTgXveq419PRQeHVa4
ad2TWzPvDtgpBFfmR08C+YZN+eUNPL7OF943YbzB+8KxnOVnXcoVIb3BAsWWsPxUMOGcpvcGPaJC
feU0ZVzd2pi6JFvB6BtfEyCp21/wyhfG3VYhC/p9hwb6ry9rwHoNw7Jbng2gIsz6CN23NJlaYPHq
Qc9OpkIPE8iyUko5bhylcDuEu6XdnxVMq/K7iwIHwwSXJ13Nzo1Xe/2mn1OQ8OoBoA9tXJmd8yoY
BI/nYqLvFGuxE4wPxBr6YccogdwnzqV4wMO35R1VrXu1M8m1xSmRWrwGpPRL90G6EZoddqkNSVl9
Ujb66H6qiOiiGyd3a/Qs893Uf3KnwvTFDziYPoKecex0F7jvlhPLaF73Kxjgg0Ao8sodYOUJvfn/
i5pf5e07uZhlMjpOyxdT96QLwSanx5P7HMIxZvqgd6fadXpTQTEHkRejWXhgSJoXUAYdedWiFbG8
EWPwrjIotzHjHWCg1UU1J5nqJzLYou7vjkoPFzpnjIJRIZQHhnMWHjZl2jvA2oP7Y+u9fScv+NeA
tKkX/i9W0SymX92npA/rdNfBFp7whTklT1qz3noX6jwHidX1e6W9CrtamYnN1vgn+BhCNw20aQhS
vziflU0fkZ9Gk1kKvEMQT8s46ZWppRJgTlwQnHej8Tz8jF7vxqDKnKcEjp3ZD0pm3GhHjWLQqOBK
U6zGcClOJYpnARCgRr1i2k0mCgeKHa9erRdwVsX6SlvODXAjcSCKDKdCtA3eJGpaq2wY7dZAqidA
DKq5D4FFx7WxSbuzCr0VGWpRK2l/T6m4tfWhKN+nGuHGg3lFn3PBHwR8nENisgV8YJ2fMgzUvLIN
8SLdr/EHnjyornFaRvxmvAWKnBL+0uRBxYlngNfx/gnUUkKGhudeRxUdhcKbWMlfTWCBo4NjpYLy
Q0WbBsj2DCKrGowWcoRvAOPzwIgTTL7G6DIjqOzYUsBUHZ+j0ve23kwdDE83lUAQbBVQ2tC7UlLO
TIP66gXjj7WgOXkeLJgAI66MsW1wQaKk9HuAv/lLny/4DpJZjs+5Jw7oixiM7q5gyJPloan3AgrE
KH83SvykBZ4OYzsa+PJkFHu86vGNzQBIjVm/gzqHR2eqeaK6w6HA1x4xM7pkaiNayIbXUtjdS0ef
6gm4jLR4124Qc3GwcRmiJ5SQtaW0yg4jLQZb9znQB5VrLJi6jv1/I2mey2ioS7zTPQE0QvyjII3h
5hSHg95CK25CSkbOrTOg2xmS8ksQELZ1/uTP8OSB6dixjezKfEAoSVL5MrwlDEu2oFOclKO9BtL9
A1xOgELqkjGOO9+3DBTSEwTgI7pvb6LScPeJWZBMO1iv7luYSllzfuiyit4/d0FfeTG1I+YYZ9mg
JN5V0twkgoLYkacvM/RJLdmUXXOAnwQ2KsQTWLizonIjf9ANhoXvXnfkbwGMokeFdD/tw423aIso
6aGLERtT3gazJDjMd+aDUcNZ+9h5e8ZX/qtWGVjyFgCPuL2e+Nz9gjGDCYuXDRYuOtAE/dZInYjE
qhLRipE3FE1JOjM1IZdh0MPEK7cgXI9fnZ26M5dJsO3nlHoT9dufZSyaIOx8j/XY2NRkHgGFoQC1
lLy6QlPrjFMBRXVhZ6rpc+zTvzf75aELnrBSalWbDC/3GwVfEwwdYYHo5Au3ABUcJ5o6YCQ7tQ7l
YHb35ikaFlC5XD3MrH2ItPHa1ojdmqMc+1XuakeLCOBmb5ta+B6tNPS2tbAFoLaeVS+m+vuGPaax
THORUuYm14IYgFciA1sgzw6Ti4eiQ0uJ1CXM0m4FJaB/hz/AsiV59ySwQbLu6kk/cPcvbmj8df96
Q+07qTUPkHZVJmaxiR8Qz3N9Z2ZjCi12F7z85gCrhvoUlmycYJ9KJwFqSJUjfjpBZ8co/6iSof5K
rQILRHtYUxP3SVriNyFZaR4ysLqzSXmG1go/Botpzc9Hwj9sNpzcc+vgaoBo3KtG5pNNY4nN9Ohd
9Tvbm0/JH/GvXC5tOSG6BUsnG4vSHZxcuUntHquUlM4oWbvoFCZxv6KFj6zS9rn78vq59RvNPG1H
z4B2O3hCSxIIevOqXY80h2A80cHqM/ozkJEkJQTuYgeVnGP0Bm/eIfXT1AucJCSOynL1JBrQGYYr
lIbdoMrw+6sTEZ59o5KsH/CzF5I0YmcKZoDfmT6EFAx6hWoav2PbGXa634GKlcAUGGUsn1L1g/zd
ncbgjSrtOemvnGN35XQvITly8G4uwwEujuvLyvYfStjAymN7yxT8KIA1+/Q3T1X2M6xkcNtSdnw5
+WOaJpCDKgQC1eapoOsg2WDxWg6H7fjclkeKpURaLPieS3LNwxxuu7lkLcNODJ/MrQMdaaLazzzz
tpw0dGibaagLMQqUN+pERnRhqIFvOAB2zYMeY7prJ6cwhAyOFPWjWaL2yYl9tkmDk3zikIJ/dAiD
dUfqXEx+hf+UaQ47P/CgHsmwU4wintSMaODUr1vmEXfI6RnzC1xiZCTuaGww9slZAT2SRdLOf1fZ
BRUeXmOl5JFQfr5E8ff7zFhoAvqv6+lqc4Ry6/dcq0XgNzrq0PD4Kp5PfiK/S3ADNEXAxogLlj2q
zDcpwaKpYj01vS562LBwNORjWbqjPQMzoL9jxdqiYMYxZIHh1Yh3ZWmAak8E5mya7WSsP1w/xDmd
3KQDehy81TFxRLrx8XrKkJ1tZ4gQ4TdO0KK/nMIqLkQ+GtMuaJbHyPsY6MOr/DS6BYv6+3s/etNM
RRa4FHB3vz8vwcLHmudwGSm57y1I4zhbQzQiheggZJdjTLF803d8jkr3acMU4X/Jhm/3XjUwGk6P
CoAI1NcS+QthWvo8kxJpU6fMHJ3Bk6E4PZMyEjEoulx0bx04lMuknTzo2lwWnsTBVj8/+tPyYwzC
OY3yucjBOWVpy4APA9typHzm/fbatVmwfhozu87MLS/RhffFRBw0RmMeHOjFDv8fElJxuBHp+OAp
6+FQueQP5Rvie4K+fYj74+9NySoDrbNk5hNvDTyGi+GFSNHZF0d+eG653boi1EF5jWqNidqtvsqy
ueHonARLsTcQOYnpVKjvsOHvj2Kb/TgEFkywGpuCBTMUliZfQGm5AT/FRAC3AJa13fU2MQaIv1Tp
UxXGd3k7iRxhEuhNCAj7o6ZubHmx2SMzrU7K7lFa1tOTJ6SVojyjpJH6urGVc9vyi3aOjk5/FnD9
gmS0Tz3vobJvnHKX2Oe4eS4dyrqtmzJskaMZrGZ89PZ0XOzS10WXQzTdHZ2WVk+jyaUp6R+Cj2sk
bL+TbRtF88OTDUBA9CaY0DjkD5s6WXvUzcIM0URBH7b84TadJjnRSpBGp2PdrbnTD3oA22Ts8190
m1yhAZ0NylW8bW3ygz+iTRuTxpW5DY6mViEf9INHfFdZ4EsowrsnAP29xM/LJGSZcaFTNYL+YuUD
zg0aPwvcsdKquUx5QlPW7aLLxu21RwNdmnREpNPUtdRBwjIcqKX1qkB98DbzqWTSiCD1x2xg8tPu
IO43N+UZfRUVn3rJ3du4gAGuR8VIR9nxrLhEkSsp4WdNsqfPz4u3oyCZqNi4D+0Y0kUBB5Tk/V2f
/FUfvToAQ9oEXB5f7tnSZh12y62veLipuqG7I7H+V+ZRPU3dbHhHazhxbfDTqt0c6bd3CtAYTXKU
5csZszcgqxfzezZvMFjrd4SjPTNAkThxTfseuMEgXI/3I4auvqkv5EMQEWrpB/Wq5b8zR98dqpau
jdLR073TVexTmK8BL2QgqWnYggKLXXnoaZatTWzy4DFxyClt0UTJR33hIOzBTls1MLLP4BSbnR30
gHUD/GA0jP0J5xDdldFWTFOvA5T7zLe8D2dNAWTRgGtzhIS/Hpg/x4tlqKB+AGEPMH6xuHD3YXpm
FzxfXveF50ZzfanzNa1JHDbJwtMgkUiVJKmdo7NrQor/xu5Idi6HiZnyPbVtEwhb1kShinYr85x5
+zVkN9LVeLVtcmMzUSPbMzTHIjcp/3kxKXPKoPWrUoe2rJhYPLx4BvnHvcTcUCym2yL+cSlioWwL
UjnY736VxuErGowAIo96m/QgZvPOdWutEyzTEdCbv3uRgg0M6HSwRFvdy4GYZdb9sTKrA/VUA9si
9IrF7pYR8nHJqLn1IIEUr7ztr0R2sibA9jSdI1QaX9wejmwDnOY2CZ8HdbRlXZfNnOzttmRqocVW
R+QYRChcEMez9rP+SBCToDvx71mK1ndVNhQIkJrPtDDB20LM6dgErx8saIgmL/BW8LLhMWFyOEV/
tEpQeUdFsaCpy9M5Y/lnqlyOXc4O+JKhqxF63PEsKYXhtaq1287fMRehv3hZ0QrhGVxcy/WYqywT
gk8Sl/BsGqrw0vJZvDlzdb3pBerWHe+bWy3FMJRaF9hAwDqY4/QPStyab249KlbD85huAVBVkXxJ
9Ye7UwjriGZ9esQBTctdeMP4XyDHVT3rmiYqHn5fAYTqVZfx9GCbb+Xk4lEi1RJvds7GZxGa7cpy
WCP+hn7+mUhI/Wi3ghsxtHycFeRSd9hGe9+v3hJVidmFjSpW41zOoC+GMnYSgCbsll4ranzOid29
QubMhVkon/45XlR6ZbREaBJT1HfY6G3O0ztdVFmo4MR1QAxlycEJlZRzDtRy2lm/XPsk4Eatzm8M
mTX1PpTZHbXpuHUyHgcEV1It2yksa/bfEpyVKHOpLCzJdcaLmd0Tury2JNwTkVoa/2KUD2mimWR8
uR+pz6498wHgHSRUS3HdjYeZBE7oy52kQz+n0AbtyvQzJxQqQLBRPBLkKpR0XkH9XawcEv9tTZra
4TIX5vcrwwelVck3hZQOf8QKxQUegySW96XB8tndt6bsTyo72jYB6NlZNVq+fyBRGeGt85HyC0wo
J34oCnC+ZV/uQar1Lbkn1KwOVM+nKpfsvGx2Es/VdzJDl7VMRHo8VQT4J3OJ3+tYD2IMDJKkuNf5
0FwzO9KA5wB4J2gat6nrMfWAVX/9dNVVA0vv8PGGFktyE6C6kpugj+Ba4N2zXEAXmjKbF3QMhI2/
WNz/jWYC4JyNwoDz7w41K7T4n/OV4CROE54K7+ZXVUZxcKZnmbvKbAKNmNgHvMEzYfxw+UF1l782
x6HjQK1ef3sQ9T+LUtUbZBIGXjnT3tSKM15sYzAbQnzMVmRPyEEw3mES/Tl0EtWPb/bOvZg8Xs1x
pMeIOngb2CE4Ka5xG3D0vDw12dSKvsJYf9iHLgZJsI+gTdk0XPkZTagGsFM456UPTBWgTrGl/5Bf
qILP9q9Inmik+cXru5jyRDMkj8AuS0KeNaac9iFeAj2RflFzevDa9qArXKeqxRve6aasF3X7mOds
HTI4VlzwBG2PtJqggNkj/ocVVSpqMdSyvAbi7Fwjug9Qhstqw+HJQaRj/rXZXsAjeLOuC/0PDU5w
tmGfiECOPelKJpb6pH0uVA5irugDJ8NFBXrn0X3U7ds4JKgJibBq3r+aDglJKYMlzqcRMJ3Xp9h5
0fZdC8tSu2wP9ecahlObYb42AhhgklY/DsLoZ+VJXqAmOAL5DAnxkdUWxbrQIStXW1nO5H9rQOTu
WgxHZR/Ix40kIyntPycRyNZvfPAuoA+bz3NEHJEECYC0B3OqhxPMDEr/YTuwK80r7BIF4KJdjfCo
7wYp43TCVmCFfnuahL3JrQ9AqfCr5Eh1Y/GorOA2AyiMWjMbIKECj5sNKiZGqrJ/VexVrSSgBK27
dLjtai8YweGrbX33gNTrQQ/8Ja/fvKQSIld/p/ZkPuslIilMvi9pFKdl+24ItkbsBjLe9zEkNIhT
+rZKmVnWHDesluiU4d8fi2BrynhL/x91STkh+m0m5cVeLPZGaPFIQp6QgvggWJds6n3ZkMF+wbeO
4nx5T3wBZfZPkq3IBUY7i/DS2eQuwzxEUz6HcVmo7v1PnZ8q/X9wM/MDJlLBwEA1pLGhRpvX1l7I
g11x1hnyW4Bag6I/QS88qgOo9OAEA9UdzUAooGUmNXvZjDy76k8e9nyKiMQe+CbNUeNLSp1+66J4
EhYd21SsEr+Wa+1gGhk9DUDGVomkK3heRF4sIP5yXzU9P+kkl7m3lN3BEWjlco65Pav91jVsjKtb
Ml99Eb5GUEW7DWgepj4IVWKfp2S2KHm5nn3BzVgvLWKD7CZUA758LRhCXRALvFXgiPiAMticfPJw
4V8pJzGPRf6qrc14VPKd8f75j6h/ZZWEaQ0kgcxLtI6NYWyILS2b1d1GLoX5lJHNMNENHfis2c36
SJtjhLMc4/CGjoMNMZokB+sqOfq03TBtagFbfKFoTn7v1TrzO2wYq7ycRNbM13ZW0JFx8qAMnvT8
JJDDzNAjasc532tSYMSTOCgqdj89PFA8cQYbhD8/PtQjbLTAK0sFCFCMbmVsy3L+wv0eeT/yTKWs
iepoh9NwhZzbaWKCkIUBK88VXyFsXOam/0MrJIPnw+OJnAVaGPPI59rL6RMF7+I37oOnZEUX928i
GCUWxDiclPUc9IjgDlapiVz0PIsfytu7sZjeTviESzeS+cyCcKJR91J4ivJa6sjfwxjTh4siuuJe
QRVIuh90XNnSzpIuoR1/8lJ0EUlkyZEpFFdxRwelyB06GbZLGzL7TUCVDssk9IGQ4BnXKj8u7yZX
lPtsEEsak7AjbetMRzZqq2h2b1VBi6JjlYs8oOFT4U1xch3T/suuKru5CIe85buM8+tWVwx9aXUj
I/NmB7qUZU/j7dj2tdWevL7DGXsn2KeIgTabPP72ZWxKtMZlBKsMUtZhXct9grKLZ9VJHuZh0z4Y
ac2pgKGrvqWLNlfGX2jZDOxADjuaJVOhZWPk/HMsFp4Nku9lsmO+yd9Ga9huTPCV4yRhhjYJ/2lh
myig4rpBH6mSqYANGo4/DnMZq9vfy61i989Ih8RvKFHYuCZZFPsyCItaxCz0dQxmC+lDL0JGJjfJ
KiwkBnT105dPAFC8j69UO8EYsuKLC6MZjcB05aZpRu6tdO0B9M41447CCVMbNUa+iV7lCXzh7OIN
Oa805g7cW8LGoyiX2FB2CGyGmESP2YhtE7k9G0v39o84iS7fm8fuJMW2ZsMcXHQ7OXMKmQRjYYzF
hKHXwqs+5NykKC8mJHcx8/Wxf7Xd+bzyfG3zfkVLiZMFAMq3O+0WAcJDHT5YyWaeVLovnQuMJD1Z
TJYwVBzAmCt2Ft+tcoh0C0fpPWZihwe3/9I1s0HxCU0UM6VOswRZ6i8SyzQ14l1WTjKe8mglVj7l
Pet8F03CQptrIXMocG2WdRKmeNIZCBpxWUO3mDk9DgHMQAZSyBAU+fKPyeo74q1eniAK4yNIbgkK
4Yawct2mMbAXto01HjvJolrshyD0Mv8atUeJIq6W++eYfBoOWgtXLOXMHB1+aPJV6oDDkl8zcui2
CuNUr+GQDf/EzmCbqNhC+fPYHNDcuRdFEza6k5fcgaQprGcKFeFWWvVPmR5EC0V77lznfGEmwRZ/
5WkCOgXgp+5wFDWgQ7a5SVaWoVQNP3Z4zjpmTHlQBJLsiiosuPMfw8eO4bJPHnLT8vk8vvBUpGmZ
4YmHvCp0jiF8cDeTuf02OeRnoqsuEm7taMQrt4IMh5w3lfxwycRvJEudJmFSwPZyoor/fPY23jrK
AdiuNxqsvH00bwRGb+xOTz9cD4WwD8DCtsV6uAINeh0V4sLzZHQR+jRzTd9rKIIxRbkaDZ4hl48L
Ie2Zo+AvDEgRh6hAjE9pd7PZjISki0zXVkxT5odaw2cLBuvE7pVkbwVNaeZCQ4IA3P6cylYzaFkU
Mx9YWxeexGXEs/WmL6ISQwFbalHI6FYL8TCTAbDZvf6MRmx5hzr2wdLmf9qdskkw+/kpswKosaru
isPsNdlCP/qkup/rJfQBcFmTV8IPW+JxbTHCdQMmlmaeTKBJxFnj9mejvY6hyUDBDD1U9A9P8/f5
SShBD6ZvGL/mUdxYBgwUzeUo7LVILTuHOWdhtqfokXtHmTZb9fSsa4EMogF8brVO+mbTSljUC/2E
PD22SP9vEKU9GlEpKf15fHOm/UWHqsWWc/VIjZWJi200PxOId01bn/5shO86ALR/iA8z2K05AWdD
GlgAdQn2/OkQUueQpv0/AfFp6am7k5Uz+/a8pkx3m+isCkvhkU5w/3sfFGVs87+ngH1PfhDdPLFZ
fYdPYWXDMea8LPtTCsc1az7Rwy11PYe4NcAHUx7baNI9kWHihAACOe6hqKCqY7LoGLdG4uA7V8zC
PLeeD5tuoyitp4lvWZvdztlfeidS1xFC9A8Owz7hfm7XgWoK5rEEhPEFsNtKw+XdpwYg0vfWM9P2
VKybyfC/o2coiELzmEMVauP0OREhV30Bky+mZc8QN1xOvEbxhHn46Tz8rNHy075+ygbzutIj3mds
NaOmdXBVcq/jSAQHFXVqFV51gICsTqx7JjZ/IvNQg94THnuWWDUX07YEGi0IrBvAwOb4m3J2Jcm6
n4alwUaYdXGsvd786XyAs61Uc0ek7GyeTgb6+RUZ4mqR+ZI4Kjpmndornege4aaTOc0TlMy0idz/
/EylNs2hrSOPRtCoFAFXJ1GVoOEM6kkHRP0DWFgqxabaQEexl5KXWkdhm+4oagID5zWXFZfMp5yW
EsHzRFqndAyQ0CbKgc5R6mtzCa7yum9D6FeyWtrEs3a7QD6DXaTl5QMPllwh4tSEwX8oykslc1XI
Zcurw8kcrNm48K1DGkDNf4+p0jMWPzk2dz92xcKUvD5k1+8tjhrplj7is/nCLBhcX+kdG7lidL01
dcEwIWj4zcZKhR6YEmGtittyRQIOJCCk7Cbbag5DbKHWxHGtdbu2Kb8n9wscdmtZndgiP+F3peWt
Nuh4YcXGZ8+8gdGE6ZBVKm2VU7Z6Y5l6tIg7+TYi2eLntdc09lFacAy1PkxMHmuZepNhGumIiuUM
rr7u563um76aTfwWt1J2XYwTNX63d7HAgncM9TCIEDjQmRy9TEy6DU9U4sORrQYncfXV0ODTlHOL
tf6q1v29TZwNRxSFqBrbmhkrcSkvKzBLxzKBur9BazlLn+Xx7mfmzyA52egVD2vBQCGsokqm23gJ
M+ZnYfm3IPVzk2EwdudcHezB23A65maZJ7nzXX4vZLE4aOZ9Ah7o08peChsJWbNAnz5zaLxxuD+o
Og7c0TM3/d9FbZBvwrlmUNm/rs+1koYBElstRjyfSQqzls5/2ZCMdHOzNpvegWqNJr/7jwoh7WRh
nslFr7U1QHUd+/mvwjTEOemkIEOlI5KscmEjIbwkQZavPMxm+bx+65JWwIXHohdMJ2K2en/iJGO5
DzetpQCnW+iQUdxZv5C6h6e+jhvlfOs4fptgY0s8jO3wtYaBkhyKa4fRniRYN7owf0iLrTsUpKwm
sbIV9WOVkUXnA1wLJn7wRygrZxFPWPzuce2izRd/+e0EHRJ/KAWBRYcRtc8fablqLpjELMbfkKvR
LEwFCEbYMPn0lTAziiC+x3f9QZify03/aKd9KilTtUhoeujZ+GfKkzx1wGaXZmcTOz47rXvm9ai4
m+aI+nmz6deqbfnUrZ0p5pGyTbXNuHSBRK8fwLS2OMI1/8PgowRMKsBRaKWNX+3roB7e3AV8on1b
jbR4RkHuXQmq4GueaDdTWq4vSZQe1/rKvYCFbhVktNSrzpRaMc7qFH1QivEfkcGgt3TDcjblacsh
Z0+6QG7QccSJFJXZOwdpAQPXO0xdvzWSxDTU23P3gtaOlVrKIkhMC7yCAaIT34EAw3mTU+qwzP4+
5cb+ZeEhJ7YXGus3bE+st/etKnZsMr/gaSKj+DdsaXM7gkfz4mq9I6bvbFFJceYHa/00/R7HmzNJ
XkbE6YuRBEsLFIkh9Jdz+KM5AzKwLsQRPPGxFk25Z4F8eVvNaEkfgiqHhzuGdAc7BFcSYmYa+4U2
H43+knM5SI2yRVwKcOjGOf8AeSXWUk6UzrZ/NtYlhIT/3tt7MEV0voEa43A7kEzLyVcnIAYntwMN
laGN6HcCC+X8vmJBicOmI9Sk5pj8N1E8FpVGxqc8ctpwlzV/K9YxLYygPMk4+zWsBY+TuKtfCCIc
3cfsWi/Ho07aiKEN/U38X4XMQaP9N0Dc5yqCsFHWq80w/tthqj11OdfXuDadAV0+dt1c8LaP3oNg
/UkQCRXk2m3cNQ3A8k8G4oIckq+KjB2MQqnj0aG9CjdoGEFyv0JWCKSaTqEal/hwUPVS5ZtJCQC9
RiRwHl3wtAoJhmrJy9h006cj1HbespEom/6TJNmrECEZtJPOcVV3B5UpVihNplsmkchxeP0U5avv
Z8qjO1Y2M6ftFsaThCMdQ6jtzvxgRN5wAR2w/THVp81vzq8jM0PgKNcCV7CTvtDNFLJHLH3BbVsv
gtPwHF+eAMAG5UTsV1n0yXO6gZmiAbHqA97OdOCWE6nZU06gbwtBI7s9wYIeQZiW1Av6ZWgMjh4B
WILGnc29a8jdDFQQP9jQNwNnnNlF9erz+DiP8SiNrzwqW26fEzUkb1DJpxKj4NL5rzcRh8AmqJIU
tmH5a6SGr4V7TTFmolm9S86kpVW+qzcihcGVtpRj40G5mjiUz92cPa3CIAJDIo2tOZWfOO7Uuba2
aPigZR/T4PELhkc+a64cxqvhsCaSgL+vSi2f63q/dEP73zhWAz1FYtvtmi5S3xh+jBa8kXUKaufF
IYFZzS9zbGj5h/1loPcHbjX4/G6nISKyUyZ4c7XwSJXkoZhYrMH/aDs4Z5Tl0NMElHRSCszBI+b2
fSajsD64MlECM5v6q0tA1Opuheg2BAd4+clPuzXoxMavRcyO4vFYZkFSKI2PJA+Sb/WQUD7AiIe2
SK2pxgCrGcsfmkPBD7EO3PA/NKzIi8okk+E16hR4xQKV1EYYqrfgtnNSyI1vA4rszJ40tvQwtjcN
a59EHKtuS9XZAE7SN4N/lEoIB1KdfrLTY9EcwshnmNxNq9ebLWeC2WCwJQEaHL7VShnbi8IIvpqf
ribduXyMhNAz14Uj1zV4QukrjnwH7yKl+Fc/bHtf3VPtt4MlDX3rKrNAdLz75soJUUH0/TpW8KjF
mLyW58aLbpUN6QghJBNli9/bnrcinQbpbPdCU7SJhxLIGSDlJkQgkA8sKLNFUjxy/tvfLdzm9TEn
VoVEpA1KWGitOivvNKN6pn3pqRUG7xbayc3k6VguyJQsaGdnttD7VW3cUKKqWo4pVSY2FUhkPR1Q
RGD/ybVfT+a/e0swRMCSZw6SsoDu/dgXjHjOnc6njDV/e6QSXGMO+nfqostJghdtE5HjTz6qELjW
r+0Y4JgXU7tZEWRIRlzfYbVz0CidIH2yTnsWHwcpZkTjrGc4T35h52mSBAZxpsDbHkSbt/EckAoS
pIflLhcZPVeXpO5iixA1cbAQLCR+BdgMZ684NZHxwYXyMpUNJZBbJKcIiNNal+SwAmxZx/xzm/vL
iW2mIcXGHT7TYlOBnDLqcABIBiE9Qk1k/95zfjzoh3xSS7RTrt4Cc2SoaEH1Jbfvv1micT8Vww92
UeGqaIaLRIdPE7lHGb0ckChB5mstnQ62SblDXMXDaEYhqJvRNbV8AM8QaLdQN2VjXjlzXAonjxey
8/EpCV3rKra8P+NNO4MLj2ISU32VGcZRWR8Baat3BfknE+sMuZFPhp2OVh10XotVwCdri149lUeU
yvsupTc9mKYm+0w/FrC47dh7yqjVOm4QKuoSzzmQyTtKvgPAi66mCvfjAgnW5S2SP1JJAnCOowGB
GI0ufdwSwHYzlkM+c/Q+gxEjERCDmiB5fpFGM9ncmdIkNlardb0u658eNh/+F8HXe+XjOIlKmmu6
n4kAkeKsNeBtBhPaCyv+HRy7WVvAyJNCWZI5bxiJCxrlnsLErJ8lVwWsTIdWu0M751caJ/5tWz6o
LPodz5LzxBKq+WzaHD3iqFc0Pv9MDcFj/mrWdYVbkiGjYbZpKrgSPqz49/TstV7OiBze1KxCClhA
93gYLBH3rpVC1UrO17mcx3sAKgj2+UkKfag63fvxx/IK8NSK/Ix32y4K2tsLlJE969XVivc/45vF
QdD0i3PpQ+XXhLn30Dw9FRo+d6vyo/Nxvvx8TOs3aueJ+Q6m35sYa3J12/EyD4MhIyDPoewey88m
+7S7MDClzNjS+6pov431fCgRs8qxCDoHP5+J0eL7/TFBe4wSR/7PnooquBr6rvidzXSRmykhgGPM
0KUvxPiO5nnCTY3Mot8ZLWNb8PAITTIoAyM87Nflg4F2Z7OoEqFHflPk4jl4T9wT8b1nxAtbR0GJ
9X/v6ZT6qzD9ButawCttACOTfvh2hLW9LHjj9cjWM/MpcyNYg7gunDaHhx+Nv3ySFg67YylbYdvE
N7PB37sScs8hHhzCqZSJc6QV5X3CpMuBNGzaXtPhYX5REDG/y0GH3o18JsQ3bmlZsq06Cj5wAvvw
2rZKqyuq16YeZpwIQqGd1hYbIvhRRdQo0zkZRwsacUyA3nl95H/uXjog395UBa30YxquBrWie789
rz0Oa1CZrXBqjlBPaPYawGxhL2JeBaSq/IRI2SdsG+GqRniQsKz3NZ2CfaR9nOdLzA/mdUFJVSst
lNE/yyli+ImmCu1m7thE/ZON7r80RoOU1Z9yGTVMp/IuC1b3H1Gg5GTDK1+wym9z4vMUVRBtgUnz
DhuiMUP0Bahw3HsB1YIri86tlaxsAGmJQ1daNf5Xv8X8V9fJUeEOcDedA6wT7sztJRtv97572ypV
J3/+96R0aVwfaOkPwjSu3raJy1UfF129FGeFwYpedlu4JEPGpQZpQibTV9ZqbHaWwOL9Aqzg3mgB
ZVmH+c4c2hL9TUxQUF1LzghaEbWOWzLtlRhglM+U1xmbN1pS4v1R5ngUyele09YlS57WA9FCjClY
1woBxsMbAdq2TQZ61M0sVWE8WYKPr25qRjSWceUEG4bXHvE89W+MHwmH2cFn6HkKb7uFkC4UeDj+
OyQaAF6wGjQZV71z9HONJsalmKF8AXhQFTjnyUsC9nkE199sWDvS7CyhOR2tptETVP639yNjDttY
eavWISqZdX30/vuimMRmyXyLQBMILApCQS3CMBYShOXlhGWMWcWAyabrCsCKoHlT43BQTRlj33dQ
CBEG5hmGSVAVeBDt7N8KV4bVpI9kmp8zkWXpVBSszS+xhuut+xLdRvKF2p6iSDzYqGdDtmeN3qfA
bCzkUBurUsXll4zRU6m5z+ThV/Ew495pMhqpRNKKlX+4NoCJQdb7MRWPaTaQNn5hYfrLqsQG+sly
wb0QpfufD8X83pRtPmAb/xAtTDf7lIs9udLplZc+Y9xUVXf4E66/f5FJDQRGgUn7QakC7mrr1IeD
dq41fixVqpnLRJC7q6gwDyulm9Uzf4c9hBdvO9EbVQh/Zexc7M9sZqHrGN31IEqIS3szNpzMh0h+
TWRFBEUuCpOEtpP17T+XKKEK2jgXiXia0MuCpA1OfhCWV5zc0AeAOAlJCvNhGUP+At/9GytioDav
92hTZbbeZeolSLvQrn7T+lf3R21HKXrXNP0/4QQt2uO5CBul1M+0I94uvGI+soIPuvkLChtUqfBg
2M/oOjF5MRoKHqWPK9mOXojVn5kDHX4nwdxigVCytQxd32B8tZng6oSfKp1dkDFnjqufHuPjmUKd
zNQfY3THlWk93eZvFRDJrNEIYFuaXwRsvGtbNcNMiPzLRYDNwHV2tdLMVRcL9g8rDSbugCQj73R3
oec2ITLv8WMA/dEasfm2gpktwXZ/oHrzMhQn88ZvBULhr1yZ/Yyc+x+iQm3Zh+c2L6xGkZdedWah
TZemNXyXvqWwWzREZZHgR/Pm8LWQZNP2aWAzSSt0CAWvUyfyoyMNx3gDcWchl1Wm08aBBCQVacdt
GsKd6hilKzGh3lQWspY6POq/NV0R3H/13VCbt/TDfgIh4GHUPbw9ARZzF2h+RILml5mUFDBwITkq
iSYdxcgQBt/JrlAWO2Dc67mTfzBkBo37+fdwfKmc+aVhOzQfxqJq7HXvR2ZzG6WCZHOUNoyO+lBh
B6UslSkErNmczvs2r/mwMJrpu7VxtQ+vasUGDoSDVk5NM/GDsEjGJQF4B1rKUZd1efUaz2eGh8MD
cfM8pEKhLzMh9k6QvZXTlfXz8+D9zCJysPR4qB/Of/hgrASy+pAe5AMTdwOH8cpXnKPX+yConYdn
m7kozLbcFD+jaN47QFyR4T5a+IDW3I+obMqCDJEutfqFOsHSYDF78T/5Zu+QU0UcaN655QcF9tE7
s3DgAhEQR3tn9IFoli8MhDkIUCARaB1LJhR6z9+GoAWft1lV0LYCNbJHQhQ9lBfn9REhUoWsu/Ev
AFsCyPqHGVvJl0GGLN2xNdyT0YRqDUlimlH4Hc2CM1xUA0zZzQpEaNBrsRF5ZbJ2YY+14F901mB8
FzBBH0t2pLFke50Xbzv0VWRbQriDth7W44/CvpplyT7wSCDhFhNR9TNRHtd6Z7CpFEhzr3Vu0s60
jMPa1N64FmF77G6KwXpDmHt8jqCns0mPGITaOJRv0z7+VWjjELQiusX+AFLqG68uQSa8X6mM8RR1
e78tz8Ub2Rwv/uujLKRPpPBS1DSEJbgZGWAPAiPyco9dhRwDR+i9W/5iMdAXpvrEO6di1YTb72J9
EP3W/7lhFXytMQHzIAnzr6wsU1knBjZ44qHH5w8dTmQGUMR9EpbkMUbNbDSjza591DKXb/VxLcMA
7KAKkkKm7FUNiO3QnG6Y2W0DbCnJfIjfGrwhSd/JfkvORSVeg+lBzIQHBybDbtXjKdCYiNeY803x
oWgs6cN6nADTxB3AN2oamxNGjqxzy1aWJoesGPNNW0qROM7V9sxmRpanrbgSbPZcENXTunJtJjer
LPsV7iY/lgX3QdtzF9Cl+2NYMGF89E4cnZ9CKEisN0yP7WIkwZZtrV+JNShTcDvY8TEZLHTy+JZE
JjzSBiSG/zhZmjhtna7lZhUncv1SGEUblZsgAOVj1G+FxfSZqL4sqdSdjJL8JVy0/rV1RlvaAYMy
uCTAjGqMPBiwAocthFC2eWqP8jRaBIDHZ2yH9bXTQWstOCZVTSNKtRfEdhpSvj17ym60rnYqA6aE
OrkVGuPE60gNTaRGWlY6QHGBpwV/gosSR/a5f9x2hE06gn28s2opNdPYghp8gU78p3Kxz/U+vFJT
GYliZMgKdqYvETcSscGWClpJSmFVDRRT1hmL3VWyjb9sPJyRvt89jwMLKBW6p6CI9lZ1hMG7XC4m
LwXHxTuYQUfmRnLQH5R9/HXoJE85r1s2T4oUlDifjbpJky15K4fynomA3pGVeNgaxIG7BMX/O4rU
/yxCyzaUZtHC5Qq/IBoUm9YnSgES7/THfxLPrioI6xBHT9PwX+MiOZ5/o1ygjS49bfcuTLVoGRcR
9LtYMYpH1oGiR1GCF3LQ0yTkTo/+U61Muc+AMWJlAhiKl631ST7Cstnb+FKmPvVCJWnz7NQPpl8z
M1kGWDyBam3KkMrfd0z8gchWazlg9bdgBrLuVI1eGFO0Qt1yJ19I793mA0aQqu0K2+FUAEwaqc2t
OwigusSPTl7XlZr36Lt5AXRGJDpox3e6XclFQMUoTtyDoI2tRnPsCZME9uU1/IYFD6jZIf/MRS/u
9fe8i7q6cVMRuVjTO9D41DYLG6pk9s3HvfmISSSDWa6+/5txqKyHES7f+cMP184WHOXDMXBQKWPM
yXxVF+86NHo1YoRyFzBFLEb21hZvLQ2auSGDioBDW+W61MxTJn9SdYRQUgMmWmpl7RcvZm1bgt57
dZu/P/4CwihelmgGjHTmTdxSCQRCygOOf8eucOHvqbQVLTBZEQv+APxGW6c80CsRcH7pdbKrNybA
avAVP3U6dFGnlVsftXv7UYy0JcV0djvR9HbclxSCs1WUGOoIoHtlABYlM8WVcY2o3GWbwPpS2YSY
xHiXZj8+aWKbGBToUq4hqwsl3538N4bSXpJRzaGDz/ggr/kSZdvl9VE4SW7fIkftjvwXJqmg/mzk
vZPtKBu145O33FwbuRmIzZy33AgYYceTFdwZ6YavTMjzDUbMuq+QHCVcY80r2QtkCmUJpYyS160Z
Gsx4TBCsaltj4ylR1oSDKWYSN3f9ojtLRTcTjfp9a0pIgCbJRE8KR8E2dLUA27cbz6u5q8YJI9TA
tqk0GQV5Hl0kzZ9uNIBuqNySvqJwue9KCvBUp7/VyhldAz3B2WYUdnLeJ3u6i/0EfjcDxT3L3TxC
7DD56SYAFQ52ghydJVDVR4SIsil8yYM4LsIuCKC391cMXwCj10Yq3pTGHsbF/y4XRtIDiP6jhAfL
uQ7aGsEAbxZ4B+eIuxPte8ZJJvVERBa8z39elX+5YbGVEsPUwPev6V8wxKStcwFObQFyHR6ZWlcc
Ls20ZdcyQpexw0hQR77ZOE1K36IbC/90pHX/QD4NJD9NOXctfo5Jrb1wsvQaySCR4qFlVHYrtan+
7cNqbEotfdvQt9eMZlZhkYDqVCfE7iVQhv4Ktph0TPWKvF5v2POjyWC1VWg/K+eu3BpXalMGq2yz
rmAKIOscRZ0iJqWm0fDuC0gb6u2OcI8uObVFXoNyoW3aCAsZKCkWeaUu6nriA/dIeD1UEUYTMmkZ
sHI3I/gYM1unmQ5nrDvXG7xw0ZX4rOzxOfSAvWHXybXytgG9GlwWqqoBfZDAsK2lal1pCZkIgLQv
CPJxG14kOcFd77TdeqiozGbr1XpVhXvfo3wXvW15qYaN2HiJJezs6esTJozS/5xrgiI6GpW1M/Jp
8rz9lWRy9SA8yeUObakR1BBfn/sJzvrIrH+MXwaKZu8pcKHilpSYXm5CzqqH15dwgQA/+gV2ReqW
kVIs3jZitUDPNSIoA5HTtU1EeyRwQn6Am53EJArcKivpsBLPFStbYMPx4EGf/KpgSlZZNQQIf9Bs
N+x1Y9dJTzyAl1GKTVwSGjpVs3YxGPSy0KthEbovyh6rKyjK6zDrI5ldsf2WEdgz2yOlfW4iGWm4
5jUCqePKRm7B8ZGeMyO5SZCd/2oQQnVHqFIjK3Ac1ysLg7LEPwtosrwOlQVt1b1FP00Tjn+c9X8y
WT5S/k7nIF9kQAHa1Z6Qax1DzB9+NTuNT9hQpQ0L9RKGpxw0Qdq2ilPvywCzuLTyeSMtT5CPEVjI
6u+hlqpopK5kVWdfcJEBskwK2/ig5SlESkTphSQw+wpev5FxBzhhEpb2FIbJikbre4r6LbsL4kCW
Y5pVCJYiihBARCr0QQ+JZmCSKK1pGK3dcEDymyaVCZbE7lDRJJ9W+cFVd9rgu3mmFFQJqSW7W4Np
5tzZ7hVzeqpVKWOxE//HNCAvllE/OjJ/vsiM2d+urC8ABdPqkYeklgXisdkQR62v4PVQaNuJfKqc
1KQuz+DzBxx8R/NikbwiLSDyDqJtE3xVoP5hxQQBsOyv2o0n6Leq7LcQJa+a8NEDtOscs695S+2D
1HVR8VoWta1N8RXN/SAv0bUcwMUs5K31FtM3c1jjzKszfjuzwtjL+6z92IzKQdcNv8LT9JefK5dr
rU4s8KHp2qmrymCS37EC7VbS99/bfUcQ+JCdTmAcNcrUXcpt0FkjCXNwgEGVfqZSCfC+6Iyl+l4W
6a1OWQ1UAZciH9Fm5Tij6mpzzUkna9G+BpQcgKD96N7eWfD9mbJw8cDOgTcrymKJy9/Qbb6U8+4w
zSQdPwJuw3wE5sUCdMooc5RrtozSLdqG+Up7zkZwzwxCTrS2eKiY39I4T1QAeTXUeMk3BgqIRELZ
cClMHXVrnFu62efW/5TJ4Y755HL3O/twmgpZt3Ythm/aOKeEhqJsRAyqZzkq2H98VSG6hVHTH6B6
gtB2U5GGia1eQW06HK7ZSusbhOKfpFBvIatNHMI5ZMcItu4WL0uI3PtQ0+eU7oNyfV0fpHKmjkuK
k2w4T59yTL0i6bc91zq4XoK3LJUQPjCSc4Fehgnje5K5qeeMRAURT8bdQrZ7QGsGWGD6u0ST/CVG
PF1BR/KVuc6bJPI5wHXRq8tuvlsrpTynkrrjMIB/l/EiA9DmdUo0lRdCM/OA+6ZfCUOIfD8/mOKi
9bIfyFzOCIjXBN+r/RIWA2DXOiauNbdauhtG+oZrsze6CfAGVuwzLZULgv6jl7ZXcJmvPd2/DtVo
oOidRVPwuzcS7kzSFwI/VtTqOOud1NKOORClLZH1Dgl3PEWmvZZOrHoey2uZb9E2Tdi/oUWaH6z+
7Xn/SmbjeAsy/WlFPgSs7f2VY4SX4+ks2j2nSysFIDJiocU8/CBORRcZ392+tVyvMdCqn6uPX62R
rQ2sIqALAmJTcCRtoPEg+fvrVluKmbYhGusTPh6tZgRiVhrxegUj+r/rtX6YSqukgONYsKKQ0Et4
zpNn5l+Xne8Y5YXi8BaVGcCDygjOhx7V2PXt2f+7NNyLGuyDkO9BMt/AtlgX76rQXRVtFgwEHZW0
P4e7tGl88squhJ69rm2+4O4qLhojhber6pxVfc/fH9Ac9lMqi1SrG3t3cQ4jxhAgEoE5KIMtCWBZ
nJMN++DMkjOJp8euOouuIXBjyVaUipsy624005ZDKUz6rCWSaCDgg+eJjdeiNPZ+LEe+qYgZzB8+
Ediibefkh9HnxbjI4tDd55f3/56TxQrmpwxAx4PEtmwmtipRNRQU9I4KCaFJqNA6ni+HYyEewFHT
f5YMDtttaBrmD05MxJJ2jKVlnbsk3CKwUpfih3T4Bi27MPv7ZvEPsgvDWfqP4lt+8gwCTFrfokZL
EwLoNLN3C6JuaDgeAx0JDncii7GfqGLHWko5XVgTViDcsUAOnsutgw4sZ1uJPtvluzBS1/Iky4HL
kQb+plBiUq9Zjg4ghCj8l1DGYJPIGyZBszb5LOzOMFvrTa8j5jaHjiGh2sZr5429Xh3bJhQ4PRFK
3TyqbyeOMytOTNPhuvl6g/dFdvHCDG+mEjvgvY3Mdm2ZeBQqD08U2sWe1GIgd4MjqWbSAVcRf/Tt
UQcH1KPUwys2EZo2P7V7cwlVwS7ONF9v1xYtDZIw+ZDTsc+SkM1rv5NGGqdIEoGEAOjScF+wticA
Fof+2xO4GrThprax69ZYRoIqd+HJ3oDNQF+flEI9FR6UmK5XZ2X1Lajoo4dIN/CdkRFLVGUAPoNY
cyPHUG9ZWnWvfM/12Ry3gylHW0HFdMingbrsrBqU6g+upVcmpvzLZBZ/4Q92ZZFeIH+AKSMfHYhX
9R6DhE+DGvbyuoORN001MeqNuLmmO6+ydcOTM6JhpYgH1KDu9/Fm2HO9hexxaPjezT5zhUZusL1c
sh++XNqT7y2eKE+TGFZrM6AKFoK8lzIJv+zuh2qBHEIX3xdibovjqi7gWzljwnJV8st2q4LKub1Q
2SWPzTBCHqKfnFRasxljiSf4ZK5xoV5S4KfV0ChPII4zq6GQ1bpkZbokHtf3BBdYcQR2fz6KDokW
Qx0HQT47s64pzEZBEN45yqPHYg/ODI/AMbNgFPi6UXSnjjvtGjYffZH0+w5vMW8z7pPRKYjAHr1H
jqVXpp4K8t1Mx0NHg4q/hSMBK7yfGaxi5MeRE2C2MfSfE0ws7IH2qoJHNbgrKCo7eHSzXwKMNuhe
dJW7DQSsPPsAVg6Zaaie7mmQ0S89op5Fo/cS9mwzo9zpKJZ37Mi+UAPY+I93/6vEwyTg8bXBSith
gUSRydSgzFxDaJ3s1/ZCGOJvl2lEqiq5uFbf0lFHtLEOEP16Jq6DtRVGiWJVMfGY3O3PnWsXE298
6uGUzCEBmEv1Dcm49Q3OQl07BgbTpRsj+z3lsvZA1tAjqWkAcjIqFUNWpWPzyqVEXfQEA6lFrAfD
kGhsW+vZ4XIjS6jLfBeV+VkIc6W7c5jTRR5vdHOHVk1Anj08Rf4LdbMSmARg55VYVQSg9GYh4MKK
DG/mnI4gIIFmFNFLt8GsUdsHStMk+OEQjqnyTOrYYe1vvGF5j9Qkk+JIuGtE/szasYFcklKgrRft
Cqt5G0Z5XecpVwaaYCl+1xH4RrwFV6VZnEMOerkWuwFwEmHZwZKP5qD6nau6gvJh5DqRb8AdRgd8
RFQlvMl00G7VvDtBAYEaamU5oq3vyjtH46i+bDdpwGousrvPtczxjoklm37ZkiYPr/4Cv7ntlJMI
vt6rkXLDvD68yKqsIYwE23XspE3N3kBWZtwBnZNIgsUcu2GI4YJlwq8/Ekx3IAx1JaoKuU+U1yi2
M7SnN5NXAGuupXslj3t8ZDLTDOIvhv2ttfjrsufUTtFWbQ60z0ovDqYWoEwqApbtJ3lgvtJWQO3x
TYbEI89l5pkUd+SEr6Qff9R3y4AeXxiCa8ZuYG57fMiplfmHTBYONNcOCSTC1+gXTkSJ94fGZTm2
jKyipHF3HERalokJwX0Ziuc1umua6Oo+qU9MQNHzw/7/mSuEgdiJlZ+brhmP1kYAOn0ERtaYk2f0
iPOLiBOJjJHRtQ/h8L7U7VgzOi/a6nIKMxZ7Ubs4unrV/JPDHJh+ruq4muMql0A3hf/y7BIWUktp
JEzC2tM1442/ngkV75UK5PNJhpnWcI6i6RqRX4nVeUW/QWMA6wIKZrqbnEa47AZWZoUpWdMiR/el
WDFkrL4VN7oHjg8/U1h31chut9gmDZdBVSKBSIi5ovAxJ/LrCNDscgLMxaVODyoLT7Cab9jYQbKX
t/AZxTE6HO3wNleAZj5VcW5SecchdlA97baU/OImFu3xTvtCAG7DAiSipBOrZyCG75IXqqc8J/Me
v4qUnPNK8W9cSFX5nMX5AYGINcfswHQRU6jQxSWBb4wMC1uNt4vutOtSwRpwuyZGoEVgVwLLmi8M
mJEJkN9guTnxkjeCVimZ/mYQuRAp5LqXCx7rQFrmRh2GcJoV83Uvj7N9evawnwfmKFAT9IsDrM/v
5eAadVnuXM7Iu12GaqZXYeUd6IqtwsRHjDdELQmu8V/e2NbKxyDNeu6Z9KSv4IhpquB3q0L26bEE
wIC22S48zIkmGsWYsYo+cyL5cBT21Kgzy+rVlrQyRQH9AhUMhSwqya89ewF3jKZtLSib26swi5hI
m9G7kvlvFVSYMHLq3jiyQ0178xqJTT+PNh3Aoh0IUC4F6VOTBOry98cksHquPOTtwhC9hA1JHBtv
gYyng2/lYP05Y6IiebMuYnT4XWXS6HzbC8Q2Wzh64+5rJtrSAgmw9Q7gOc6Chsr4m2rwBC1VWb1q
uCfVxzw3RKFOBoAKc3blZeCUn30ILgkbkJMtW9UGfPJslZtumHJu+QTrrofWv79cvg3co4+pZCKc
1Isqjp7LIp0dRfJKy6b1lGQD6Y+2y6LM0TIwM3L8sm2ha13I5UJ/rZW22jmOnGTmaxDQzvRkTIdY
yho4BJ2Ife2ktAmIU/5x61L6GAmfhljDRG9Fc0mDfxfaX4JDWizExEvsC3DS9sXvbSztsrUgKiTm
8OYFN8YaGp7reNzQjJZattaN9t1YB7CNuJMvC1gvB7uLL27e/ZeKbt/uio+W8sOf1L58cJuGPjtm
Hv2sbQutIIRy6uwhCc/ZxED0Fws1dTe9o9nzvIEnoV8o3vf9NAcjHCvuwhx8QlzCWSNQZZJjOUwk
PJUU9e8mK+UjnPy+AdIHLVyidc2h/5TOw/Mewta5f+NyUBwqUVNw8rWhpPQKWW7dliZApGGmx1Bs
tvPfF5TjI84Yei1p6p/JWAZPQcc4QdT0H/BwLTVbi1JALy1T9zsh6CJlhGUzvkfOkiT0hHEDmrJF
i4CkC9pG+ceGbCINqNtm5Rj3tTM/197rn9vzdIctD1WTkA6/RutFvrxR6jrXFbgxQmQxojARoNEc
AYYvHk8VfokBUqeJbUlE4ZqeMrg+x0W2dud9DbOhMhQvEYCA3XXG7e1O91I/xFBnlW2uTB6aM1WH
hfy8NjAJrLFpJq7obRJJF2BzLShIW6ovGuZQquPV+tvXsSkpUog9iPV/vnAkV+bEFKKPkWWJ3iH5
mZSFIu7YFKIUDdgPYFM6glL0z74nx4eL2VMAMRJx8qA4h1Gu1QvckQ1pTzmAcBq5eyKWkGIfDG0Q
LlMmDLXWUmt672VaBoHr5CKeJZ6SiZaGEOjHQDytkzHVic+ijHCipf9fwvic6Lj3kG2bxhIIpQFN
UocKsfl+m9oGoZ2fv0PYYS5vDRHOAjay3kUnykzAY4FqFkKF6J/IwX+2YRFl88l3pggqreX551R/
IQQ1UyTtkZjaa6CaW8gy+4lr7gzYljK32QpbWxFlHKjw7fQA7MmoIfaQelIOiuYFCdvM8cK1GHTy
ES5X9ZhQzfrGxoD3uS/rrxn4Ue1PZPgA/xTON+m+NPMPdT0+eFtt2VGM9Ww00vtcruu+b9hMf0Iv
ScghGg3FNDZBPRZkArJXZBp4h6wK2xKxZTtrAsSVOrAm+SIKQwoxbOABjW+zIhakYI0xdQAgxrkX
ew3YTEIw3UFhsT+9/QRsarMaja3UV2HnZe1tugL1gjmgfS6WAb8z0sqp6DTXwVLy2LFlTQxaaQli
QlY4GT6uA7MnCD2DD9DbLR+TKV9Xi7Cd7PKf6ZBCCz3KTYdNeORM5bJyO9YTOQsXU+kBCwFVw1xY
2h8uhdl4cc8wW7vQQtBcpJI28gdKgJ5QNioolNXDBJCVZzZpZxDYk4nfE49uBrsaGBTE3z3FSWVX
ns1NGp0eVw2+fSCFoaDa4Lppq2VslFL1bTuTZ9Id6uVXxlRproVZJvNcS+pMZ1s0+OfL9l8YLht0
TLoeEokFMR4RP6qUTYG+96snFrSx47GvvoNk6s2W1YT1D9gLGGMDKvezVJ8H1DMuQ/7Tq+NKmGOY
JD+K67IUgRpF4VTu00v0ArnE7HH8BLAIujwsXABG7iKLKvIH5ksEObsFLzS5DLwWFVQo9U3qlZqc
vL9SD5Jhddr7si8EEhUeIa4FFEuMVjbW9xJjY7RQ7/MbotacZ4n5Ipvy5v03WFCDDqR0nqqLhElN
spiGeBjQNAL9AcMjGrr2Y6xLgY0utcqvn0nTjUMbhlArfbjAkCMlVuIs3rbzAVDpC+zKnPqlTz4N
8FHHQlRGsdgQuJe4jJ0jftIjiZayCKlrmxIURXzSn4x1G2TsL8GAsbScs0w3T6GThk93vxKfwRgZ
pNwSNIKkM+W5giTA3NU+F2RGQCwSs6qQZiOwyncqq/z7mqMhNMaz4uosSe05/uwyjr0p/2Wldg6x
3zAFIWTtJsAu0w9iFy0UjHuxNpsp7L8zOEHMJXPKOgnnFM9Jew24DazylKBMWRc7AC2F/LlcRNPU
8Q3imKPJYug2mxS+kvgHfV1XgArl/TNb2ZCPYUhaVsFsdy6sw12dwyq0EM8b3Bu4vCpZCh2totbb
7r7G8Pt8Ie67+3Aq82WEmxFymLwSOw+xHgj97lGFuml8WpO9Rne8MM7k+Sbhw5n/Hmnt28M10va3
+QUMf91W0PkBsNSlZ5fWDykbrNCmmP5MqBhS3WGVOrPqyWgvZdoSIBnstsexZIQKHNKlkW31yr0T
MmpqOAZ0sB7Ll9Hu58DWBJDe36ZLOaJoYwoIL1MijGzySQLPePZsUCfkQjythDzYcKCSeFo5EmUo
sHafTxLjPQILU1WkYl3VyOGkPH1f5qWtAjh3OI6I4frzklwc7at+EVri/02hHovGHp/kycliWVT1
zfreuF0kyw9nIDTgYamuM0y7FSvlCic+iaD1jVSKzSu7vP2EN8PD06mFxWbH94MhB2pmo7dRk7B/
9EJdf40ss5bnOgKc06dlweR3/QuvbGUg+lX3wq55rfgPapvnLrOKHykfADE2Ole9fH+CoeISML6J
mVhU2NDAJ/YSfxaSDcE80Cr2vGjiJAs0UFQvHlGK5yajn7HV7qjuwldDHRy8pE99xGAKXTA6bvu1
aM+y0kEMh5XeSSRrJ+eIB9PRd1U+KWKzLpOW8cwWuyiZvGMuG5Fs2/m2usAWslpkRVxMn2vejztk
vPHymQSt1+/jQAnCdicz0JwKW+joZq0OgXKE4utnHpZg/m7jgC52k9q7vmjXmjMuFly9Hs5U6bOY
0wOBRxGbqK+SLy90xhhlP1U+STOibLO0wlWCCXAgA4GjptO+jRkajg+FpvbsiPWVZoOc7gv1msm6
n6i1r/zaVAM3FwyaejBhLOkFmhy+Tw+CkZt8GlzUcmmoUryWEOlrvdZQS5SumBVzaENKe7xTy3t2
pcK/93d3+yi9gePVMhBKdcoS5Hcr1mMuib+PoqciJu6VSBFiP+9o2oy9zrOHdQuL/40RNSFN8MzC
fsfJoEvcxeMsqr+czV8iYNBqs3Me2eHT5w92q2T6y7Zta+7hwQQ2FaIemztRi7+18b41jFI2iTx0
hCF4rc6nrQzzgcOiKAbMKO91CR74/xllUtoEoa9LKRQlTHUzwNTqN33dBQkaJYbdiYyP5TW/ldiv
REMwTB161z7vnG7m5VPuKk6sZAnkJQyYYi5pvvBR2o9gowwRPSmBad9gHS93rBE5IpS4rlL4u0jN
+c7LnHCgb26QFpvbO7pv6YhAyM5i8lFmN9KoAyeZ4KG4Sp7GYI/hy2ZBmUe10y2kq/F/0nx0FiUR
kTiMABVzlKXiCNUeknbSHGNFv7rJNXD6TTgbCLfdaZLxf+m5391NGD1QkqlCtUp8j9AjmSYeltCn
yqpYegSOqPO2khW1eHSm0LJ7QiIkmnJMzOhKjCMhM8vfzH46ss6rrJRw5lAvgZH9mfT8+19NWlZk
9KN9CAjqJc9tOKkmb/pPl1GRmFyKU3sMeKEDVghEUqSSGiise1nvzSXmWrw2sAj0UwdvyFxkEltE
p6TMk4ohMjTUPkb2fkVhozwE/IDPSciXTfMospoLVCVUd+jQRRpIs8wKUu7BoiHeWsI+RPG9KeXk
R0TJT6R0QcApIAY2ywo3vuY4pfcDvwf+09ouggaa4dDuv+JDPT9bdguN0k736WbhaU6nLNmCjiug
ZUvaca0/+83hUdh/P+FxfY1bQErFPxAhuZi0mEgDmR6C5ZF2ZJcVl8GlHWUPIF44vK5L0DZg1K2z
yhV2hQOxQESz3ji2fimMiiBkFncrS2UMdDzxZDKfr3Z6E8a73LhcL2cAXReGt+hgTOPTYyHjwq1u
omFtbQMD3qgCI3UGXTX+6vj1iGWOMbbPb5os/0XiQpqasW631Zk94Ll2SM1DDEXousWdtrEKESTl
lKrzVRgwt3FnX2bOeo3FDF2q9xwHifjVU0XDsqqQ/sFwNO3wdPgGU7zfiShnXDudZN6e+Hfm0Y3Z
G/4csxE/Y6yJtQhQCgjaJMipdZgBL4JhXF0VW8kwMMqyuGRx56wkufdOP4jBnrLTkdQ+RCH5iMao
PZAnvVnFH0xPcoEMJzaNlMPM/a6eSJtmtvCKdYyFNX7SHGYtjAI7kK6nKH57qFHpEv3YcD9f2+om
XI7VwzYMyYOVpO1f4A2G3HFbs4tcaoXR56u2Q3xULyilyK0QXczdPUrhGa8lcSLu+VpCVG0xwn47
vyJHAhqZQlm0jXpVn5IfSNgeEumhWEsxcgAUU7Uib/MoF8CwLJLFWH34KtVhcdzRhU9yW0xcchn9
igRn1OlFf6XQgessd/E7Wrw/VhmYoH6XMhEy3pAx4MZ4v7Xdz4Gi7hzfif3KjhHXLtm1/auNOkTe
uRDimKpSp9y/WbiS111EDpYK42uVgxtN7RhOcfQO9tAGy7ze9ICRmnjrUeSpCh51fKI3nbdEyUH8
tR4jVWOQ7epWUpJuyLh7FInhrFvFLD3celosHP69gb6hGWEB6VKPPtGA3kqUMf36YSMm+fIrbtRk
Ia1TFKgp6mePBEKrrXBEk4s8GdrWmWc8imIrQVdNKn0Je2rx/nj67z1yXY9Tkj5+wWmYxIHxnDpO
C2mPVprhwYMpU1/68UW/YhqgDSjZCzZqz/qybnLqIatuhQFwSNTWi8J9r0PQ2Xj5i8u0PuP4MRlY
nnn1DX5wwGqQ2oh6stOn25Rz9ioIm7+RCfuWmSQIvIBx79doCjPqeiWIunJJfFRlWzNRxZ/FCqLY
OciZJf5QhGo6yfwrx/5o8h4uT8TqUIe9jsI/rUpUlapkb+cFi6xCP+uB0YxxabsurmPCCMBPno1m
l415AhYv8b9eQsMnZYWZCQJzHklU4ZiESmkkIqznI1sSmnlrIDhzelRhYw31T42mvvQbmE6rtmDo
+JUoNew4lGgZx+wd2YNZsKpAk0Lr4dLR7kju8JvssQRL8JXUfuZhm7a/h6ifnHC/e2c/0SCWjiob
EOxy8p+IUuPA4O1xUOkWp+qbjZgKO5iG61EVh1JnMC32QOCinmHWm6cxXRkvMaiqXUXYjbgodpyA
c7WET1kCIOTaAGofgsRdmymRTBTmHQ7VnguyWhgV6oPEs3ayPKWvdd5qgba7sY5AKGCCyQKdLg8A
gJVwhyQVutgiT41bAj9/sNn8yozcsaVA4hL5KqN9uzMvk+b/r6PMmIMU4We5q97LPGzU6di0Zdg7
zJ9S38yrjhm8Avh3q3pjgHdb9pSh5D4bn9hQ0YXytZFEDkrzFrkw4ovENK3u/NIFrlANkY9XAWk9
M3QGExf0/xTTNqTaAjpyWHugptCZ9AZVt6xKl5xUSQju6s1UfkvtmA9DR/1vpjU4vTk198Kgs5a9
ANcyXM/E1Kg2NtTpZiuDy+sy3KcurrJrhTRR5aiNq+jZJ31osZXcULd7mZoTXnJ3OFjnA8zH89hx
C9Sz6CixSC36OttPnxsrk4kJveS+Kixfr3SHd0FRiRyvBMuNrh4GcZ4VeuU/cAAlCtvJgXUW09ks
YXlwjmIyzd7QKgtnpuJ8HwrMRedawFR5+5/DV+EF4GZR4dzVqHS9EqnXJFAZdkXGnC4UVkq8vuE6
nZj2bKzcLkW7UOiX/wqLgkEI17YQSepy8dqdIZoYOgs83i+o0xGzQYEbBDw9k3IyP+dvldKXpKK2
ORSpS/0XQSxe7V/ROHI6O71OMmutEnCgRPXJvgg9bVG1RlAQCyPTx4SARd350NmfJOMqgHNKw6Vf
vipPlmy32V39rO59DvbUPjgV05e9RrYhTHYd7MoemPEJAEpswBGYW6QWbWxD+LOI9olyn2zE6z7u
4jBtnzEw6K8NeKWkbvbayvlscY2dONxA5PSaFAiCWjy30t/cttRw9ELJj705dTELGk+8fQdmGHqs
OgOGc8fptCc8GW9vBVzMZ+HapMKcf+ME/5oqaiY87oynqBmYUYl/C9bHbkcNKErLy49E3Pw67PrD
j8I7ymjnJ30PbPmNOGb9iLCxN7KJ1anYi5NGRwjcZiWn7bM9WcxcLwTDiCPGWpToiQtZRs+NleyR
w6UjGxhfENRINjOzPlXhMMGtMeBjNcippvDOAZQBCj37YNcpKO1TiiUCT9jFp9JjGGfScMzJKoH9
gEyAdfjyK2bWr5jKwltY6+ezC7qlqxZ7Kr7tYRWjqsaHXujWchW1iacHfTjqgBARnWb33H5v3uka
H/DFcfdWDZWXRAEJhvmCzguzpVhsetOXij7Zr7gTGuVtUZuW+xDU7X6ANkvRAYhfHYBDXons/Uke
7IcrZ0ixlOQlCExJatxVw4n6+bIGGFoagbzatCkcBsaYTYcYi9ke0P6SdrJtbTHrwdtVSu9aVwjk
i8+ArzDF8x1GJwNpfyejO3TsU9j+1IcwVLQC06lSIhOkCU9b4VV5zLHjSwrDr8AMyy2ZGmDhMAQg
nSFDzuTYHXAZQPf3rNIofVQYR4/J0C2nUmsxPtfGF2R59HGWyk+wfw8PkIoo7ai/hLJV8OcKs4qM
v751EHobHAIrNxgoY/MQuNmgKJ11RpLg4mAQzbNNu0upeP+zYi7hqlDGoC+czrk3fWOmUDFGaK8z
/o7jE2u5oM8takys2gUKWrpTbRu2p9eXzzPKn2+dPukXGX+yMPxLuzvwxMc/HSVqCMOQa/FjDEFT
gfsBsq+hRGGhs68Eibo0E6hv9peDABRo20O+bTNlFs474bFkyp0sWJJmssNxclrqLpCjptg5SkEY
kBFgB7K/YKamT/rlQdYoUew/lWUmwReqzDwwPi2pq6fYSkKspYRx9+cG9kqAgaja5JV4Kom9AW2X
sVC6o77GOI4hTGiClqKzDz8tno1jHAG2VYytnOi/U8KXp50JW+m61QyETRh+B2o32wvxXaY6zRks
+o+PUmUPsWOfCYpUmQ7ONxYZq0sGQPS2wWbmdDDpXSK+iElvGOFjqNNMI9mUD5ZUza03dWWdXixU
oPQzhNfihdYtnkhajDUxt6gSIhxILBzH6Qr+g+cfsintpl4tRWq7yPQud412w7V2HuGdYo1KTfVG
uKxsQAISatWKzrbFRVjrm43yuTp2RJtKZLRGJ0ZCtkbwwmK3rIV8eO57hFR6EIxEktG6CVs/GQkm
fPnx4KwYPu86bGHlFHUnv++kiczAK9mSajPYKN7vHCL2x+R5vovgfJplISNKRAU9UBXTsaW0XkGg
G/r65aecCUm+s4O8CPH2gDuouisWD1/qDdzeKoRKvAph1s+N7akz6WaCE4u8Zn0xTwqaBJGF9Zqq
kUtcAjSpl2vpKqQVIcQIJkVK7bBZVzNzCuB6cfR3IwQHe3vohgmGW9nn0ETFR8sYF5ENuAIqsOG3
LCCJZKa3oPthn4TAK6w4O9PzQLOA/4uPBwl+dvuuKD0G3U/4tpAtvAJUt3THy7D3+ZFnZPENAN5C
Fc3QrnM7mxo6w0lMdUne8Oa7Gi/7bE/CQfKiNQW8Zm2JUvufffcOvDWYD5PBMkpxSYtM7c8mziIK
iuQgfaPovrNbVvnkA9c53PaRtuEDAfjcxQyGa6BCYmJzkkYNvYtfNv3iOqRhrKBSo+XJvNGd0IRV
vH1iuB42cnjE/Y1MQqLjAlP4BmjWDBRGeqkenZNgAQ9ARK5ppgNyAfj7Vj9ttA0C2ZkOstF0aBnG
rvEudI8a5/2q7JZX1mq+B6ghUAtIeIG6bPtWGH2pR5i00uucXJlwPGulqDwakTGL3BPszcEm+Mle
JKSAT3vjpPEld2S8hqm2ZXgPkrLyTs+NSkXerqE5tXjjsoaMQEb6hodKON1mDc6CCcjjCtkvk6TC
Pt81c8bq8V6Cyb7hrDgwnRwd5IieSfdM2NvG/uAE0F/q0lq/3nLDp8lfaeD4+HL9HGTtFCspeS5X
E68GJnkjsv+FwsJiPqgKxOCnabb1vbeDP+lws8zYz/qKBdWRUss3n0cFxyy5sq+Z3YH5tJqMH0kg
+PntphpNPAXkwqPjSuJUEqzqXexL6OGpuWQOrthaKtPFkG7FrTHLN2/NBtxXf8QpycJN8onVfRLq
mtJLjhBNMVe1wIdMJn96MoMfQrS2hAiA9IzLznCTithMAzrhAuWJ8OpVIaBvm9prFhAz6k4jUMWJ
huSjQsxiTT9c/kV103shnqCh+mGHyCCeUPr2hDtcGlWNCk0WmrA86Yed6OZCfi4FcJxAyjU3uJJu
OwSPy2PqjdrW9y1z4I71Dkuw0E4dqhCatSRwtabFY/q5BZtJa0ybjL0Dx8qMUkeDQ/OuLvwtO4Sp
Ey4c6sm8o2DvnRlwXR7XobIhwJ1VfNo+Qn5ITQybQ4TMMU5bymszGFtTQ3mwYzfclQP9pNRuKBYd
aTs9WkhjJH/EuP53ClDtC/YvYrRCrVhaNaeZWT8sE1v/Rb39KP0NwbdKqtZypA3xQMkAnrxYOJS7
M7KuKwh/WhioWQFfn94/t8my1R9YZX5HlVgCtiW/5aZRK0JOmLQt2s6W+dnZQCgxa467M8iy7aW3
+Ug3WD9k/e3r57pmVfzxlxdFF4dgHg6LSJq3vllXqjxYKFNTyonrT5id25I2+7IO+FE//qrikbKX
X/QLTEiGO+tG+2bhwc4AHtcGIsEK2+hptZXMGbn1kbRhD77x6YkgVdJaCkanaMr3OkhrhjG1BdlO
WzytEU0pc+6CJnYrRU3I1AjqPI4P1s2vKewfRYBEEY0ly0OmXXRQ5dr8vbHVDN5qj177qUT9Y8c8
RYeEwPGJgZ1tPtSulWwO4ftkkGNtbMvly1C7gJyCAT9MA+3o825zerLx1yV/ECFdrX4ZXAcl5GKc
rma95j1ffsGVRtb1KhUAmxzPbtjVFJr6Nnruek6+qlx7iYd1zsZ7bwwI7ODASyPGII78RLjLobwa
aqFzFmYBpzO7qZ0WRsEhK7Cpqo8fG+kE7n2YfjmQn0noGHWlUVss9EmwUB8NNN9XonI7FrlE9Ymh
Y+HFv2lulP+oUctR8UtM6K0fvurmQAS7cig6pBB3I9QdD751gsoUPoY24XYKMKbjmm4YJuCgqNXe
mS+Jdw3IFpQXgvME9nuF0QCWuvuqc/QFMlKnCcpaI62ndDusYyfUZQSmTWp2lPhGrugO12gS4lTm
IG0SXw3WtYo60DTvugs3Ps7PoU/bQEiP53bLX12YfrV2cxzhdHOADam394FN4/eoBL+xNj086mHl
jb09DTZ8ZiIKIxTBVCOBj4ag+Wz2agW1ntFSmHxecEbQ6K4lZ5JB5jaLr9sNOdMdKjv31qNjnSY9
WdlEpEQsJJ/tn+UXuwvlw0QOO0z3Mj0HY8lw6KrZxrgz1cyOod+E4Tp+iUR9GkutpU5788QuUs/V
MjBWax8IMQDXmW7CKoy/0//qf1NxEQ2i4alf27GdQhwgWHtxtsN3Dnr0CxCNgZx6L8MHA+3XhqFk
NLpMg76TDqRo+23W15AlZQHUoVhPnrM1c85KZy3skIMtv43khAOm4rstUCtuJzIaH7Ai1VFGBn/b
dDJ/0bqkFgnA2O8g+m9J5+qA+QWQ/X2nkI+zdRbGqn1pa8amOf6f0O/MBA8y1iw7GZHHZVdX//LK
JvcvQF5o48Vzu1ficCQZlyyaJOADIn1oIQBILKM5zyJ1XqRdhY4oGNZVdyzQfeG7OLL0xiN/jy9i
iYW/MPKs4TgL5BvSw7eOvCm240kOpFdO7y0gaG4fKprTsOaYkhz68DEGYbFjq3/2ctjBcH+bupz3
kpZ3EoUftmzQCNVxwuF+pIfapRbelYU5fs5QqofUStBD6W+p7+MbwFCp7+qAdO1VYUvmqH4k5XFa
JnNAdfLxBZDF2zQj5wolqhb/ijWKBFE7xOq8Cferidy5dbtlfd+SJrXNg+3uHyGHomTfTOjY5c0D
5xmcarhO4RwfgwIU8smkv94KcnZK7M2LqN1qq+NMAFOuNfcFZnAuhXd/LgNHAPF5dCZXuJPgXzy6
xbqBZgQQQOedmrh0vtigbkHGShmzckrbtrULaKMP3D6G5wrJXUFQAVcp1pb47tuwM1nvJiJXGzLo
qr/fBsOSqeiD2Ip7I/csd+G9LiJUQ5RP+MbrZLRRPRQtH5qWxnntzCFJ+qtKEUniO+1S2P7Fz//1
w3cWU2X7Wd3ffhLNvW0RYmE9IKqmvGdosaSd0ri5XZ2CQZvqyIYgiVVgVYh2Jph+dFUgs8N1cKKB
MVC5omthpSQxLufn1ZQzJXeTyDgq4JMl/xtyIKyJ1Qs41kRztt/XyJjr6m0gOzaZBt4/SnR/wZlb
0O59ihUg+gbE+0fb9lVV8r1fya4Po3+ltv/B/0XeZwgh6sA3iHWvGeGSfJ6wTh4dmGVu1z69yeFb
ZzNwLJM2hG0iweCh9u0zjydXy6r2gKZQda8wZzaXEiT769cM97+q62FgYxJ6+dX+Vrxulx7RMynK
YJUyuPUbV8LHIr3OK8oaoBMGsIsZv2zrE+uH6ZfRVIVoN6rA9Tl8P6xoI5p52hA7jC6oQeM1sVgO
X/wgL3eYwT1Ip87ZUjfgK9ktFD8EFNnHVxO4R5oCt6s6DQARmc4sNkNIWQic9RLI9OgQo5zhpmqd
0z8I4hM6RpyG6A63DXFLIKsDtDI94Ne2dyH2A+WgId42rlg0MyltfVZmvkLtzqvAHFnffkCTCaN/
rqdyH5381gDpNk2fejoJ1JoW4tKifunbgHCC4CL+db3qfjKtWqoOOBmA4v5M6SF+EK0Yxc+pvytu
fnBQVnN+tE+XvJb2sc0ojA64pp7d6kWhGf7Qi6UwaDHQSh4VrrpZdPnGrZYF57c4ZSeUP9rKJcvW
+HmvMi8DKcMJXl+lNKp4m72PVeaB7jn0f/n3teLPjKoC6BPtHkP2B9Tn7jrrsrfkIYlGa0M4oGsq
ybCVLDt3/jNTPuMQXFEBKQSr3mK7p0Hooq/lIVx8OEqonDUQdMGRlV/uGBxWlsOfMC/GTr96TCJA
c2zbNAuzL+fEqJjVMTKHYs+Rus9EXremBo+tCDyQrzD+pH5Ck7p7kD1g3dysIzczc8225/nX2qq3
qRbRezqxUzWyk6ZjGiUs5a/3KxBlTs8ZtqEOKbOAns1e9YY/roHign9ndmo2YiRCKelxObmxEbJI
HzugCQ0XAwzHL0TPxj+1WltCECtEXzEFWpe/VVqYxP/4JAD9yrl0ngqNvsLjL0R94V57Xh1xZo7v
ToLaDvcCEamCq+z/oKL/3Id6xq+x1StUAZNkh+nZul9aku/z0Fs/AcqMuRH8AhdHAiT4gYOeeNiL
/YAIk8QXP/6odLBklIEsWAX+p/gqeLCiycnKlRKynxt9Gb3t9eS3sAb/82woz/QEw0BwaflC65BH
SquTneGuBzyNwRV6bhh1pJDRnaJSlGiI5VWkcVwRXJsR5evEEZ4PLxpqfu9GaRCIwb/T4r9zpvuF
7YJAeIm1yPD+FH8NGVfoN5mWQzFS2geuticrUZ6aoUll2pmWh1AdFHJymf9uAGpO9ZY1OdcAhCDM
4ysCH5SQxu+xmHoiB3z0L74KZxe9Dq4nRbCibcoAHpf97EoaPBtK18I92jkyPQZDXxsOKCUkZ8Pp
tC9ZtJ4x1yttAq0QRi3Dll3kqU8WiEqeRJ/Tijh3G6ZZde75VoyxXVh1DqGMdkTq5kkLAwIJPK0B
Lnaqs4o8X7h2ni5YbPasdijMtPJ6qy2+pEh9ygLFD8ya23iokOQXfHmF3BfoLYge9Li4baFNYNWb
U1GX1V4LttYAsUdpiTvn6AgV8l8Wgu0gp5dpSRUVJaQsXf1K+YYx2BjYos926e2KIoMGgoILAJ/R
tjbfXXTVfeFYKDZiz4Ua9xPft8NXWTRsj+cNxx1HDpLxPuBBUQok2P6Iqv9cWIQX4SHEBDS0rlew
CVnTdHOMg2Jc6BZvg0wCZWbP0IMfndpxE3ka9bVZBubihOfHTjK7owCVUJbCUjpCwwHqKwlL5eTy
Z1uJMPYM/poYjk0QAuH18F4H0k9o64rWCpWNVOA5IwT/ozfF7lS40HRzmfrYPd/HztKPPIYj1XVR
QxPPE9Hwqgl5wLEGMjAG9r9IhGuqtNDmZzFJYo6rkicD+CA6ITzbVsl/z4NOtIlWVHoOvZmlEdX1
sd4+Tyx23jjPDcuORWh5kF/lIUvrBdFdWnLdC2Lytua86hojj753DyplwiU+o0UYo9NDp5D5nrmy
vK8MPoHb3HIIwUzHDKF3xiSZH5RzQaDM7C4Fg7tQPHqdhU8ULadFpkPJSRqnS+CQmuqpfrSQ0ZtC
jYux0A4VEUqvU3qvh9fdmFIn9V5QokTtZc8C7FrHsLcgFxp1lHEOzAJmpRgXg6lB5G9VuyfhI96I
unutcVGYM5oWgA5EancxG6oBhhOhF/KOhYmHQAOqqae+oS/5FIxxpYryQY9fZ6pREyyM9Yx9RN/X
vj+zSRyVYsNzEK4a794XvX9OY3Smmrzm6IDZNPXZJUyXcBE9c3rllZR80ToznV/5jPdmHoy6bZF+
uEfNfFcgFT6JPKQwJIXl1XN77cQcfw+l41Lax0tRn0E2z2QMwmp+C31O9GqXfeY2PfERcWPFNvYx
yXWLJO7lDtexqVfABYHp6wqeieq6l/sUp97Bx68ALNkbnIhJwF94MrogHZXZU016eHHXNynr+WoX
LZ9kc22ah5z+LBPoeE3LClNiEtl28Z5tTVNeqLs0jJkz9VUkCdTM7az1BZZeVaoXnCLQI2Ku4wjM
gvM9Cp8OhT5ERihI7hlwdq2qAOi4r8uApWh6FvLNqlyx0BWAfeZxY8vFYz+x6iiuyt8bpj/FkAEX
BXxsabvOZ0NUfl4OrPh5vzCl1DwpaZghs618GaaUSnxhRN+PvkeFvdfDdQvEMLajtw3fBQj96EQ4
HfHUg4Zdej3Im8ji4imZV4WWTz6h3Uus8IA38nknx4h9l4hC7nKsNEL/B3NAByIBypk+ji6pjQw4
HQsC5t4/qrBk0E5KYvk2AemQAhKNXnujIttJu3eKTatXXqxR1HKjKWy+yroAA4FAl6fVsfbuZupH
gOEMwscEWWl/3coMuC0uU8k3KLhqPjuweNuVi7+3JS1iYMLk0Qc6fAOLkxEDQsuX/XFcxV0ueshH
it8cE7lAjw1ehVJAmWM+Q+I8FLD1+3GI8FBGnr806becXTK7pXvXHZxjE/I3NVOUPQqaCWt1Bezw
X3O+UkhBYp1t9DkUfZXNSk0bqLIlHg5nFivtZcQN7QmxU90hJK2qjCcZId3QNFoYleMdIm/+INug
NveRt3kDlxpjXuQzJlCwoLYSacwiVBxFBTkblnfm7/m5Ul/tRTue3KXdmMpX3lzNkHVrwEOLiSnp
nBgxt7UOEwM4VbtPZz3/6YYIUHc4uSNHcQINb2tuoA9+THlpbfn1mOmdIoPtt+ahGAbBbtK8pNef
IRe2DBsG8NeNzAjpkbhkt5DkaVFp43ufmquJGpVfl8I8eFhwB/2l4V3lGVITiwyP5KKIrOhYdeWc
6Zs3GuN2zSUOAnwkvYCVTBi+K8l1txFlD09xjle8b47E1hopXdoB4Vogb/+/Ud3Z/ZBG+tkvmE7P
rv58OZlw0l08Rd3tQ+mmpmGu3miHScGsb/TrouUp3BHcKvNsftWFXaoyGycMxic8LTkLzsO4wUsh
NZ64pPlSrnU4PjVOwdN4H1TlKvQBQe4lsmXGgN7LQ33wk2ukM6LQ09iKdT1oYr7r86FpeYqYZO7P
nOwhQCSqxckqebNjRJhX1L/I08QBTcr9S8roJNRcAI7VWsQlOR5ECNFB7Ynn1QI2dYReY0cotPiJ
ULiVCMSBgM9WpTdTc8HLsJivI/cGNvOvlcoM73zC1NknYxvSOjW/RKWKhqyHoW1bA4uaN3Lclabk
acI6/pp7jXg82hXEhr60ISncU1QDayM9dyd/bnm7Ap/zkGOmfCJ8or3O30jXqnou3W8XN0VXfLXw
Sq+1QExD9E1UqGpMLTsW+XJiYAroOWkY2hTq0ndIxJu1p3VTB6YM7/jTukmoHw0bMzPGYccKi5/s
wxI+qtLg9Y2sBYsbnxox2RxMWPyq5OIaq+zpSfS1QWbxVFeYGZkI6mIvxrdO6QbYLIPJ1TCeKS9W
0CDowMk2o+XKiMSSDDn9u/dgy6RAm0ocL2fDpsqcCB/JIPl7jloIEAIhn1sBOlmoq9LxQZyauokA
ApqQp5q656FY4didKwjjH9qYm4gFDCW0SjUYrTdohxmgO41YhbA8ea47dlbvtfaAk1P43jhDmr9Q
4PM1zvIcAbCi7a8e0WbOmNvyrwJiQruvZAqUp6nO0VvaKA6wqavbc5ANet6I6ZRX2RfPdGKFWVY5
8H95rAiMDZjxyE5Fp/zsH97lP2IjgONWvDJKrRDWQzJdjwudcinZJRq3PW3gofzlGO1VD2HuikJJ
u7kFvDX5dPvBIytdJ69287ldw180db3rmQ4cbwJYpsRerEbV8g8TufkgXBMMmTQBHE323MqVVciQ
N9JG7JBTyWc+zx0Yv7ATn5iz43T+SZItbul17qY5uq79/oM+zG2KNeEq9bXndTXXmImRRMLlJMZa
zO1VXUgxOaTsLSt/Jbp5fajVHuVlsu6Gk0SJHvofS9kuwLwuEe/8iomFg5T4+RpjdnfHQ9MIKy0U
VzDttGF1f9rxMMg+cGJyb7mXkDvOy+JYhNKfgCzvYKad2taFkx6rRo893SDyreLYfVFyD2Z+AI8S
4dPjowRMfVKNgifGRvizqyvuKjxDo1O84ksA0YyIH/bVjkFO/6qT+9lQqRTw2dTvBYYiE5LjOoOu
8qZp63ROVrStZE4G+JVOvB9ADSjVreDy8Pmn2C9s1+wOYCYgsEYuIdS7eGapLnmHh2uUzYuUZxC2
yXyGasqHVNIpe48/rZhHjo5VF2XteCOIwwFv5Bu8w9nE0tjWjOBMSIIPGU9e/mdg3mwxqL80qLCx
ySdFOgdklvv0i/0bGgG612RVizde3OOW2XG7HLbk3j9XoBPb3awH09qC7/4JpUH9pqHseJ+ccx5T
xNTjRbRm/Ou53mdfwUtrZrjFRA7BHn+X+Qge6xzqITHHdxYBCGtodIUdiswHnIgmNZUjDNvKNq5g
73+To1WPsiW91IQkinLjSjXHFI6zgA8pDZuMZ7vMVzITwu6zn9/M34/mNi58UxagrxUIbqwhLCFa
UcMfw1bYDErf77HOhMejgVyqKIRQIbCbxVkkOivHhsmMCa72C3G/9lc444SER4tJzaxFrR0NAoVW
5sSTX2+GuszPSm7nTIDXPWMmAAfXYI6HftlryMIZ3yCOSfvpbhGbxiDEeObZ7Ed9n9LH+U5vH/Wa
aSp8Y8pxEU2gJuCUHIkZs/7sVgA3E/QbF0foBPQohKoYO7hsdsAT0enI4UQfjMcDrUJ2/VhJXnQJ
p5z/5O0JTl+4MWPjieReh5NayvVCnLqgzi/xBfVOabVvaDFNYlrf7YHmXv8kdoC8lZaDEtShQujV
EswWuUvFQ1A6J9yyayO6JTxoQTQQFUigJrhrRVEIcz54p+jbpKx86GqbpEpZYRjjQ8+2myziVecG
Ev2TV03q4lM/lRNe4XzukL+c5dAj0JtjH0W7Kr1mRYyOl1yx5Qh+ggcm5yfiWTKn5/svPIOi6j5b
YRdxJKAhTDCUksU0Hl07mEt3x2IceWmjeQwUAXDlwq3a6pL4tugrAGJVPE/+ESI6GV9K1QcbAxkD
D5Ir3Qk2EYn7OAp5nIH5s0irntIdHhSkDAx8CtiGLdbDTOwH6B5TI7KjpzgV4x8AkFCHSwamuloA
qXbOrEDqH8fNjn5Km9PZeys5mthhb0N4unCx0Ti4cCjpH1oxvHmbTeRms1UQzI4AHn6Z6ClHARqp
5kaQOvwXUlA6qI/3MSmCecHyC2+ZSaqgMJ1D51H1KfyBVbZJfxQnt5Q2+Eg8vmmKv89V2SgPFAS6
JS9O7CCFXCraNS8crNDJrgcb6/Bq9mw1zoACTGCpIISKXkDqqS6U54ZEv57VqWC+mGwFtnB0l+V1
fzqrbgj4KPxkSSLgkf3dzRrRIH6KlA83kI91GgaWq7gYMJ/lYwe6MQONMR2nF6GVDuzAx+klua4F
T/EcGjgVTb6MT4cMJM5wTzbipXTxm5bOVRm3lTx3Bm0vbMe/tA1jCc2rvXXHje22WS4EHtigxxZQ
9wXzLMFInkzw6yu9Aqyjfiy114YFg3uX4VVgHuyCB0FjzhHVXX7EHkMvKZ7WZKxJbolKEIA6bRXR
wQ94l27oVN6+rcdJ3CAtMP15L7laUogcEHTRdufNQm8zhGm2ajt0iUcS/TOxs3Gny9E85CXeBC+t
om9g68W1hWukEkW5XiIujPNCvky8cNTsfoU7A4B/aevI8MzU5o3f+5Pjfkg9lLaGnn7DF2sHJN0H
AsZikOBD6s+OUpKZ4Z+kdI9omtR7FINlvDnhdbJAgP/XoqBcHQOKpTmOhA9FMcJJmr0lbB6XA3iN
NrIVzGJ5TvhHb3yVLIRDuhY9OcUuiIN1MbueFPRvxilLuje2nGtYQtre5dY2jWlJtB9dfAs6HEs8
7t/VXCf9OReDMON7qJ7LJhcGT9Qs3iEK271Qrx3f2HE6xhzrLp3gS4LmaqCNmUV0JsNh9nHOjwSZ
BAr8Yj4b2WnOUs04IsITulnvNos05hKpWb00CiTs1Tte6zeRTfm78YRgboaQ5wFNq/x4jOGu6cqD
Bpk+kDBSiAVqgYc5n3YD3pRd01MLmHjW4cF31cV6aecRKI1evgp6XIffGsevrZCIgqShv9/rGNbI
woJ0CGy8YXtoQWGPdEjVclH8r7/0FqUf/OmDHquB7iqiEmn5Wb3ulwUGmk6hHRmqC5YUWwPLg7l4
+MuMLBEgcv809aYQ+t+OkzIQ21XibiDKqapdbF8HX2HJBWSjV6PUU2lcf6kCgbYtvYQ5ISZdOmms
oGwRBkMRb3UElVnQAtkjaw+7AS1xchCtLbHp+hqa35pCCMVdcFhqW9IFrl9iwvw5+8dA8svhC/eP
pOzxu2mfCUHoUykYmvxd9+bUNo4vMMqVKz/Jqy/rerjhZnea43p7zwMtTvGKHJ4fFOmPJfZcqmNx
HMHBWj1/qRPElpu7y6/2AX/sDLqZDyxp8vIx4mlLYeaqRUgIiMShJbDTBbcQtBmwemd2JToIPwN1
ThYLlamHqWdOQRGwh+36Y4ZiWGNGA7ROgxyeafyDVbnYIGr+jtMGhhR9wladcRrJ20QtFsTMj2PH
GH0x1sDLvbasIpSrd9X+FkFtWDIzxFCIMEKqy0CIsx+r+TC+l7u8OIP91xWs7iprkEykraZ/qZ/6
Z4GFWXGGJ/uJUrW9QLKBMgUnzm//bC3ZBLgBNK4u9r/hPZ/kjYfZDSfrcAhsnu6U+XoTrvjmd/Y7
0/p9mnNc3gRNf9ZjEtYOE5l6P8fIUFUcO0jEh7a/Qhutr7ssEOFRUm/ORtk4lLpRgGOOqI61x+z0
JtrMXYnGT5B5ZfywGB6xZ3OeJk1k35+2UYBxkyUoDGZmCBY4P7IUTl2mnj1xoCWlDsIfClWoNv5C
XI6UNIjvExLx5GNqDxuuVKt90NMsHEvHLpjwq4/WikoxWmHgZZ55+InR1oRVR94y+5Qa+9/ACwAY
D7vS9oF1mcMTkVbWXmj7RC1BSDdxJSrQoXAg/4Z8q+kv6+8R+2z6bC6g2GxqTSPbGV7IhaUZEHIz
1WXDgD7zXPgVQ6DMCRhIXPzwuGvguBGEtVE7SydLYIeqSQZWyGjZ/5TvtpjS+UkWKqr//fR3RxM+
jC39MenQWR2MkDSvgVD/wBWMq+j23gqkciT8xyBPc2KPVm7skRIeSnE+g8QCppfXI+7cHyN7t7jM
6OHPbfgYV1mxFCjkXJzw47jtz4N3iHDXxHCFMt62bl+CnSkFCByLJKzt1IO4BFk7gLqwlOvdHvW/
zMrodwyqhbPJZr9LZvDxywk1HZxMKxCi2cU849d73fImLHvXTtjGF5/Oqt/PDEGF82Ukc36ODSMu
qREFOIBD6vqu/A2wssYe/FN23J/29wjx2RDHT2UsjAIvXRlsdDgdaXtXlOGw+vqfU3iN/RGj6p7K
zjVUFvkisddzOEau0wDcXPHMIb+a43u1owCfIQz1OjEGXV+x9eqU+66UVQ2t/KkuSkauk2v7fYy+
HXy6ZaBULkG/I3PDgPQ0VBBmZr5HsOJkka2WtHkqxiw8PflEIoJ9Uv6lefaVkXN5MTl2qiXEU17G
Nu5VpK8ldwAgLWp9z4jW6QSC1z3ujNRUY0Ift1XBSXlXBDM5i9cv0Dnt3WvUkccX1LPfaVB5yl1t
DEMLqafetpM94ygamAkCfR6Lj4/nNyeNUEx9gLf6CcEuLmRxGvOAutld1Ez0yd5rquUbOOAByN7/
0r/HgpGDoL5qUTZtyKQlMuMXwia9mHJXJPs4tiFRsOm8SWFSY2KhkpNQ7q5V5cTFX53VpP4S38Ma
QDDGGHujhXvumeWt7IgS9jh2JxQb8REf3cLQ5EfaMm9auQ6U9gSApGHf+55JnspzxrCObBToMDuf
hMpZFiycx9KtoOXXufbHsTXiTY7pWOlQIKi+bfuEv17yDyoE1XRqeTwzbzc9a1nhHWgJ7KnHi8Ij
Lm9Fuxs3S/TGAN1NkeKZVHh1DyKBIenz8D+hf2sN7iKIVgY5pMXisZglWa7k3Hpxj05gN89NwcmU
Ira+2nGxPyxJnrOEk3y+L4vmVz8Ba/hP3sYzNycz28TjcFXxxxjRwI1QgC6Ik5Pqm7RE76bVpD32
wKUqUVFg7yllNUG2XTriUDZN2I2mjw8A0h/DOYbotqxVh1IsdiY7sq2vEFRrxQSkeJ4ljPdych4P
8NUSPCj23UyjFx1NaJwlJeDYQtOL4ZXLpr6z3GejGKzQ2Iuy3aAdIEjTp2vS+k1z8utrJDeNe6uK
pHfEHpQNateLmJ5kBoKcwAKOl6czIgmN3hO4jamoOoDTiCUMIK328pNRRX2szAidVPoZzMr1fdcT
sUvNuB7w6OFIlyTgfhaRkgRan3kce+/mYn5oZxUZWgvqBYjx4ntJe4wT9Tn24YdDjhTvGLhj72yh
a5OcKOrCN28ENQJzvRkRI5gIw1XraW/jB40fnqjhiRfkIlZ0gz4qE9PNsbaakLfaccysF/Z7E9u9
J4jdpJapqVDbcaFx2fc420YHzMFkIQ4LwAn38uXlz/FOmnW+TiQwqe2hLXaeFtnsW4th4nAQnr11
V4havia4HQFTngPj96GIMG5VJgNqkZCOyxG8gyZBRzGKpXXRdpKOkBvrlj6KeuJmqswln+DALYUu
8r7YAOAGjzNdvqap8C5hLQwPo5nGQQ8G2Z0t7NRoXIPlSsmzKAxR+IHOvmAnMtijBvKQvlM4Olw6
pYM/vHfszEOLwafSLwdS3CAr1pNxTDA/ZNg3gF+EhoyEBrjts0+seK9mZGCCaxU3s9BWZPY3RPZM
9Exi39CD+pHKqZ7uSpqZqxTl9ydLCAO1HyJ5EoMa0hIkkXqwj8aDGDIwqZ6iCTj6s2ivw/nJsKWq
0LLqK1m+Uqwc2heSB2J3CK7kS9rqWr6Cd++MtUo//K7uO+WB9+10HtyL8WII+KteZSeDt9atBbv2
WAVOeLfkDwIkR9oaG1rZuv+LYRo1z/VYgo+DLf3iFZoAeQ+5N5KNAe2ds6X00mmQPF1BQ7cSWeMW
d7AGS2QpRQhvASXw5sAsHvjBOszeTAvwXh7WaDHf5qRT3gmNYy7nBCM6u7EYElcODpBPaDdWH7/C
94XsLN0zXduipdgoM6hQ0jpfaJRTMXjWObJNe0GgaejwcznLS5n/xl0SMwkZvTloxm6VmDvUyqVv
szt/2d50Ui+g1rfkNiXXxWSct1zGZNZNdpZLoXCo6yvxIcpsMloaxDdZg457mbpWpLwniZh+YRWm
5feBai/qV/9nxI7nXnxVGeqej+3lZ/SAP9t32p0uTWHOLshdkVPltau/pRmx4BHw+tbu3ll3olqK
oyzlozJ1d3oZv0WHVEazzdVQc7kL21SKSoNSSvixvobNLdA0Y56ocT95kaoZd9WEMQ13e3Zd83kK
e1eWZ1RxswLzFSKO1VKKI1KCpjwFptqWmHBfTl/Ntrx0dc63PC2Y4L8Acct66vhBpG53iUWD6x4q
tV2tBaV1OYcG87YcFQy1WAJmNTjW3ACnjKMBbbcKZ6yacwR3oaB1q8DIFB+HoZbiM1LGcrFPblXt
PlD2Igxoirvi5sT48F8i6+U35UJjt2r/t2XE5dJtfEJEnpdEoVYFPMyaZSsO8c6+CL5qLWARq/J2
YrN07FXgpFvw65RlrUc3hpdpiH0Dfl6odVQZbNyM5mw01wAl09LOV011dJuqYUi/DLOEY3ylLWZC
mOZjC5O4y2yIOP9IzlSikWxfWMlvW3htKQoGf2ZvocxEmmZF3VWHOPRpdzCkm/PidtuNJ2a0zBST
UV74yMJ62PLbMwnQzhYL1rvkHY4QQL904u62iU09RhjV9bVR4ZC3d3Nm9/ffU0KX5t6ZcwSpOgaN
nTxy0/jrpJA+PmFABRlo9xNto7otRHiB4OaWL1vCLuTbT9247wIu7U2QGs0frgiwaDq0UkTRebN1
gbGCBzN5fAjiHcPcHgalMM7muFvoyf6Yp3BcZg+aMjpMhp9QtH7rSQZ1QAN4OW5aGbk8rhxKQHDb
GRgirziwdvy+rnFgM0BUvzg9+4e7bEeTfXm17mWgI+GGWXPJeVwAhbPBcHQhFS+NWvp7k6F/fXOD
k9LwkgC72Nq2Rcydt/eiZr/2sCeWoweVB++lvmpftgJSmaVt8duIoSC8/IYzfjwrmF+lThKaaM2P
ayyNSkB0KzI2M0LQNDKqGirlv9QOcrNEBHO92PA9ORuil25Zo/XwpGLR7Em/EzwNGaThc/nvV0D3
Dn0yWvA/xvk+6suYITrcbi/3BbvuOwculFEb5V5//WOiGxfxZ62tj8+ZFqN3gJdHuOY27Hzapglp
xx97wqUqGmn1vfyHWgkAiwoH1/6NOfl/LQM72ZWDrEENCGfP2Javkc/o3EAATwoDoc8tanEFbjln
ChGSZXcXvnUKSRQMtC0rMEWSvVC4GEBaeuekwx+YhPvF2QrXeiMFmzy8sXS9qwdnpOCtz/b9IaI5
f0LqhSQpstG/Xw8LzYuqXhJ9CHEIXQ7z/pAxScF8NUSIY6EDO8ftRABmbNplBBj8cNqd4eRJhodA
xnAfVG/Jxsz/DHzQYLVdTE9ynWpq539p33/ow8Zg3x6/9GH8LT83EWJpnQtbFxZswgnDUd0v/gxd
4XyfXbclj+/sXKcjvwl1fy6XXioXY1oCSlj/2v/00BeSlMPxXgLEP5iitHLPnMthD1XQljpKVxjM
AzwfI7SuZSjv9BvM/nUKar3NpxWRGttCVzXP2VbA3/9lN+ON50GwtfcaFJ3oFmDQC6AcYjKQNvDd
XEnYR9MeL1OdUA+yIot6Qy8wMH9IR3UU2I7PLostegdnD8fO8vmPegYtmXf9L45mzq6Ea0sZ4/AV
Nan5uv1+QhcCvn0qAmbLNQg7x39gNu5ecZs9BTB8+D/TjnhgRumRAmu1Yl72d/JuIwQvWBk7AAkX
VN0yebYSiOnWs1HCRW1N8XWsibHl1TJaIlpY9LzBZbcAMeJjdwcXVrfDKIifvYmRXbPZVWmzvST+
bWEcb1pYteobUUYwSKM5WolX8v/sR+VGRjdA56Jj1xTuxExcdK00SuIjLYrJYdszL7jYWfDUnvpJ
+pQKaaAnqfCKgoMwihHeEVu9LQt3MwyiyyTllCOd9x/Sq4K0AuxM1ClyxajHut46/ZOpb86h/JpT
S6QLZhDRlRLqa9+0bP6DHoti5ranWUilNqanPYBXX5e6sf7V52wYrqUILVnaIlpbdprJn48vozVk
vV7JEVfkR5WydURLuerdAqhY/SHnane0wGlaVWJ6R9B5/3x8syRFjmQFrTvkzMk9vG7swN3p40dg
lErZmwk/qcO/mkREhgZBVwhcB5BF2z6a1QNQYrsQPbp2XwKtFXp+pyMVHHQEGMdsHdVGr1x/7m9r
/KCE672tun6yNbgVC+bZ2NyLcW0P1mQo64nCuhbVCEW076W5Y9bzGqgJlJ9w5JL/GvOKYt71NZ88
Xfn8ycEXWjP+eWRLyOwT+wgYhvRbqdrnv7xz1nB2rMItETTkFqlCZpwywMc7LMUR5oRGVKGF9o+z
FBHYgYMrZR0T3jvpwOFKHHcPSLJ64f31c9KfNGOvdssnpfehH2uO9ch6nQ5uiRxDZHteykpCALZR
u2bB3B0Jx9psgA8hc5HDIf4v3VpUn4YdJNXDyAtTtgLBNR4YDpc/GemZroWQqC+PDVtwp5eDg26y
8nR2NT1WOA/OtaD2Fx6M52xmY6seyJbO5Jh6IoSiURJFd702lAnHhxbVpyBMuLNkPKbuCwb4Snqo
H6qR8sZ0aiA9zpchhlCDwFZwZWG4rKDZq8OS4TjkFXEIq1aEEZJKxdD527/WiosRXfOAnhjbassG
XzpiP7gS83WOIueKMEOqubdYKr69xGhjBQT2iHptGR2NY+t10ebYTxcYoHyFZJv6FIz7tK9qoGiO
sZjW2QRAXZU+MyisdYHOW03zod5KMaHMjqsmB4fUBJFa6SKBmnE7Il0Ec4I2aEXfnybyb7tV2CeV
GMEn2dnVsXJ2Wx2cox7cBlf1Hv2RmQgdj4AH6sHtg42LuEELidcs4lzNUEkHjLXfO4aG2/Lx3qaH
WmC/n3Q+6C0dbWm50aPRvUusJLENu65yuf97ub6VnjSMRV7313C/w8n3cI+A70VKA7YNDv0Qa5oX
zYqqD3Fc92kMJHxTkWASqUa2/sPFOhwGwPw8CSPy8nRDhLPh9vDd3eFiQpnl3B/mUnIX2RYhIdGp
BOufgHcB5kuhzwiLnLoUNIjFBr7nUUkxQmh7KjyZDMqLK1VvmjSodQXWhi8VxUmvCBwqD51X+OEn
PBczCHMaX5z8EFp/bes3yxlDeL6nOH4uX29uTK6LuzbHntluCzZ7cZIOP8YyxABrFGYGTDOhM40g
VDo5EFU+7SjvAHaOt5PKq4YhL0YchlFyqwleyUP4c/6Muk4h/V8gHsHiRGaot6vecKhs0UepnLDu
p7xld5i6JwR0HWL8AU0LIldtZ3r93iT7e8labCeXhXeVXOkJNVnnQDUweVaZN7N+YGlPilrTJ4Sl
JGQTEFz3p2WNSCldvE8E73WvN3bMDWjTxaoNyGSqqY08WrIfjepKk4c78Z3sd28z7CkMWiuVfC8D
Lxp3te2WIqR1JjJG0eVEdZ3S6Zg49wRfSyQQvb6RNiCCY/X7pSGT1J7tLXjSLwEh58+0Gxt1drby
UBCGU4zsp2vGZsiPxQXiLaZh2ZoYXco8VfI4o4HkjcnLheF8TLYjFZr/lG3tgwqRY7I6qHq3ctDj
7czPaliMJuiV3OMKqJDurbo1faqG8eQORve4rTjj5PJMX+8/6sk11Udqm87PythjpKPxyGHzVvri
+v+tuMuZQPOHxJMksLcsZC1ZZaRmT2/mv9WmUITlH4LngfKaKwwSzXvaQHELd76KjOMAhzn6wdHw
yZYxzesuVTvRMbM8UiUt+xqr6mUVjShwoK1arSee/B89sw7Ob17Cs4fMGu9pjTTJaDrCLwjDUAtG
g2uh2R2/gZvuc2sKNKLFaQr0bJdA7cXhahcrwza5WztdDhManjJ83Msxyy2yhZ+b7T6ioBxCsS16
ytH+kOOHQKPVxf26iUPe//M2SYLUjxn4a2Icg22Co81TV0sAwZKf6fqsflhFnBN2ymDTuXn9g6+b
AxYXsfpYHTg64EpeJjbQPiif/Y2BakoMY6sVIO/XHUBe0JxWi4+R75Kx59sIydK8oOdDzcRiPTNA
T3cDj35OXLJ1H4z3DmDzOZaNeo2uyhSIPwr8N7vP/uyJ+3L3EbgojyZ1jnS4LXNBPUEI3SYEENze
WIDDdOBe2jzlG4nL9mnjVHHDKUGSKyMBvTOhx82aYIdMwtVIQwVgcpj5PQvQ19ZlBiRbxW8j+C0n
R/xD+USa++J5XYF53D6LwBwuNCQbaayvGWujvLzzYIT3jEAhjxpMaCxIyIcFzU4EiFXo3J2a2QRn
PAhiRzF+0M49vaWIDnYyMa6NqD0sjKLathNZQ35hj8AmJvclqna+w8iafuR9IRq+OnFrK9XxQbtR
78ohUFJ1nrj/QQKM5f5b8vManE0XiZDis3H4/WpodSH0gifE4hUgP+eMcFsb5szDRLYndzznnIHu
hgwJ84e6aZem1vgBFdqPx+KR/CVXQP/69iCfHIjuTvnBKGlVOdHRnOaR96flrYyM8sF7EfNa9zRi
QI8VMCJyf8ZEtF5S+2mZVj9Zd8mRIMib9QLMLX6yucLjq6t3vsbBtbtuyQR1ZxusngZ0kZTk5t8n
M5mwQxLZsQXUuOS8HxwRjP26WpvQdNB7MqQ1yPNTaw6/hmL0aK5N1t83EMBJcEMFtJwX0Krvq6vw
RX9/dAPzVdJEK5/XtI+2R2kE6vb9+EaQU4eEyW44cmu1l1ugvHjHRZiCVMXKllXgsIQKGG6wkrAX
Ulnsj96ZvP/aeAgfY1U4uvm/bYOT1IRieAMZ9Ra0EhbvrtuFT0tjZ2mB8/E4GBQ+KHarm9gi3GEJ
wp4aS+Bhw66v83+lQl94PPA0BaGnIDLr/PyFFAVwU8SWbQtJhhQgn1j34qgXo3kUHFjB96blmLvu
/cWTydoT8Gk8cRVc2gwyQBROShSbpsrXqRByfxsPAlDHdBaIWkY9S4Cm+ud1L+YfbLcnAVlCSHH3
XTPSwf5F/xHvNwnLw1+CutlrphN77K4uaIQ8PQdCI1HeXPtGAH7SBZk++V7NzSD99arskqUY6NDi
8lL++DSJMBAEUO8Jym7Z4w579niBpJtUNC2MpwErHuO2On3cPnoq70LKl6FYDdUXVI092N3q+f62
kxHEJBdV7B1c8toFp91CFbKv1hVmBpHlxoKqj2w3VSflfttggXTW6NL6DDXmn99FSC01l59e7HdE
WCPkBW0lHbXCItMS3uc3eNVeeBRt0m97XpfCn/VPIZPd5y+3su/RxYTzsTAKMqDTdC518vgb9H8E
E13YBp9l9wdmGRd2CjgyYPPjzguZkSIBQYYcBodXtLHlhnlt+Iqfe2+zjQdoG+zMImzUgVoV2FmB
48hoA23Bk8/dk2orAVr+GJyLI0TDTkzekZay9OZT06HDUy86IziCMwPcTYG55TCv+vWRV5Dkvupa
V5nRIuwis8kIHfSjf0gIm8D/3Cw4OFfdlYm9GzlQhBo6xUgW6bKlWJ6JZlYEfumLScOFozlZy9tH
MbwWecl0dw6i7I2gmbOyYnghVHkQOgIv1arhafPbCPLvgZSYate3sLliZgJrKW3K0GNUL8N1X0io
xlpc9ztjUJKOiVxsuh50gp6mXb9FR/1klbR7Z3Mu6R8CKsACH9A3ZaHsFiIsxz0RMe0gaU+adMNy
9CFhmBCznPYznfnq2xatsPmFYnDC2AAU6Zxh8FPfFpZ+l59jywYFUI4+wOLQ4lfDdcy/ROpeM/35
+hyTWRgtzoetoNtJJtn/XB0sUP4w2ChUC+Qkx2QwivF0zutBapLVUiwnF372+2gq7bBKyi2uJgQI
u7w8EoY6n11hx3jgqpcoziwapHFnioFFBRrKNt8M523CVdBz4kzPBWLvh2EZ/hdg2DV9eXeN3/95
zIWJ71L6ofgeNSiH6vGVDJ+b0BzEDc1FhZ3BRcsXsvQZJQY89yA9W3dOQwLFENUzbs6dAh+X5NrP
dqCG9r6OzMCsPY/8HOQaz4lAi9j/Unj19G9wv1LsnE59hjax8KZ2k6zi7iMwgMKJ3Uaevia0Zc6j
3Z8VC6woIPfevdb4yF93WMMBPcqSfOgIC0I6wEOYBE1DmPJ+Z4gOF2riH+UJDSbGP6B8URV7FAw+
9K5kloR7+K7vboemsKRYdyi1/4U5JN2omStIeNkJNA/io672Q+Ko/WinuobiVK3pjUfQEn/T1JYU
ryinOrR0z2cKHXIhmQnMU/4mvsI+rqHY3gjERq3Lcp0uwGhYo8mFky6U6kvuzKfw2UIm2RPFMVIa
umRZFA833D/SzFhwd7X+Gjok05FV/fSgiNKcg6GXy/ZaleYhOL704ov3NJBK8caMgujzyZvss9XE
VE3WmwzcCsFOgoYy3F2pzz+5ff284uPR7B76jrmitFIzAtD0S9JdUbj98hjbEaZMtU8HYE4XZ+GX
yUOS5rHFIOC1/KEhHSGrIPuXPY0rYsBuMda24s1Zf/lu1oGOqZ+7ttyrRrpiURBWVWMFlMiPMosw
t0HNIOfTzqPiDpwAbqsierRKBiCxT7PGeC9BYJ8EJRGbdAyRNEDzbHFr+3dfqFBoUqO6midKMQos
2DdDbGlQD+diM0AotDxGvf+aiy8yIMk2z9XnHtyTjOz2MvmTuLTwk9F/v8r4/sszT0hYW2GS11Tc
zfLMfLRXL1iM9+XdwjjJnHoHanBA8Syp7e6K3F6zFHmjnaokfZIabK8glNMQKlOey0yZ/NPBDw9I
LfgL67FvHzouwGue2jYF8NDcwHoNn2nmqG2wxw6gqGOazSkE84BSOdIZe1epdZhTHmSnN4zkoQmU
eWdVNXQGI4uNeDSgBZn8JQQv9UBTdQpdrcB6ytV+sHYQgevreSXeYDQbMwtTFWt7VPmD5wytdEq6
abP/bAQY/Yj9GN4U2pg+AucMzSPWg0YUIIXlyfzrT+esDj7KqDQG/xk0nSijnmLvai4JYlOi9Jyh
U6XE9cWcJb8G6GlpFyTuS5lWjj6u9Ld4cBH5pzxZ1H0OiiOysTZS9BUJWojTwkdW/Ts/ocsWpTEC
I8AIRnToeqPx4TowSEGv4yd1bDJoG6cZDlUetoESM74MTmP4VKCgGkZbLV26ubbO6wDJ7QX2wDJ4
Z5YQ6sgeWMt6xb+eU5OTkqE/8bIs7HLccUnSEV5qMepjnBlOF/lxjsOxo+Bzuvi+J01eQxGWc3d2
FuajfXnzx2mVITYzwBFNii4isaduOSHNCZERmyOe30Us7J6aAAz2q+sRt6LlPCnoAQuZqepQNdg3
ojaxjCHlYlt7X8aAqu7b1dS0AiRoEYPcR3li2tULJxnJveEu26sFuLTIRhlMucnBSj+NpBu4q12l
Sd3BBFsK/oC5JpgUX6WzgniOi/rqCo2/p8/8e3ELumy3gT6xdDiyycprCB8OmVwKyQh7Ty5tw1J2
qHX+0AQTM2gWaGwV774qPhDq+nq6/EoKn9hfnrQ0AgEeXyeMcKoR1D7HX159Qihs31JqA0IKPNLt
Jj4vGxTgAh3YsKOJRGbgCBV4aa+KSYV6yvAx744tl3qBDodJGsHGA8fv0jygXYoHFHkqXMtyLBnh
wWLXNuLe/9UcKGxjl0IIT8o4i7F1BQsqt8aepJqWvx+RnQUbyAroH92WiHWb++AX7xSdFpJ5Lqgg
iYmEX8KSDbQQpZfYaz6Z6eas1b0EfbL+L88XR9D/aCn87Vr6w/S8vtyjLn848r3Fn4VvggbWxHFY
UXd6mwQGt2XA3YO/qNXAhfZSwEsVt4Pe1vpd+LPEywz8ZBWwTksgFjEA5ST+D8VDy2gkCdUj2wZC
DjsQ/o3yfOaitN2vOEZugYSwiF1tjaHPZ3dKuhPcCcyg8EK1ojz5vVhiOwf3W7BAy5qC9BhY9XS8
IAYUNj7G02ZXfPOHcUOuyAH4FePHoa1OyiGmaGVHf67M9bzQtwnr5Axlj4BwRfiQuETZM5a0If1F
Wi0u9vcvsW32eSkSjwV7cUzRisHgJNE7K8PfRV+FR8gr2jp6Gl7AbBZFfDRG2YsoPujnCbJEzBZm
FzS3nT8UQFcso4oSslIBpA3xLfVj44j+5IBd+KWm9zyl8h6NuTKngjveZk/LBpnhfJrYzA6kjqWb
jEvtEVzoZk+ovYl6UYGjbQmVhzSl1UX3Qa6dkrB9pQULvqz/OxUSuKs9/kV/Y+V/sORGjLigVepw
2sHMEntlkeSVs0pDjl5KGJok595rUFg6sYDtpZ68JKLiPZcv4wU/+lXnBosYzW/Jryr0/5wxQ2x+
MyUWyEehVxoMEZ18P8ckxZC1fYU2oTGFisV/paPoV9EuAgm75tB/1TrODUKdZalNdb5IFEBNefmt
a3VmTnmxTiv2mjsTi1ruOkUUsmJcBVjKNkuBrTIQTE3tMn4W2DBx8+iEFWU5JWFTF40hOrLSG0Nb
HYwP9jlIZdke+0CGXx97W/hI+IdquAAtkbaZg9Ie9BvaTowwXB3bYxAXz9fW2G7sHR6/9idn8jzU
vsP5VToIY+XB+xHByRqIeiT38wy3yUwhBGt6ZbfEui23aqEoS2wS6oP3CKZ7smRJfM/ydcwlxWce
TY6LCpmYi32SNqlTOcRJEQGp+S+woMPcLm59ntqVXPcTt965Yf3HkMQ76PKwemISaRED2nw6/3g/
RxC+zfK7fOnGhAWsBbOoM3sbO66aFAPHAf5ysicJaw52h5KGIUhxydWDNqpGnuYWrR4oxEpKg+op
o5G+Bje9hISZSgpfE6X3bcYoE2gomuqbvMxboN2czmIlV4qDKPkId2VHioU/zkYE/QtqpQ0buZj5
uAZ5aekZp462uxEt+ABK8+Oxp00MSsPwQk1G7Mu614AWHEH43lxkFgBZJ8jN8NDFOjMGXREQZ5ur
eI8am9+wyUzxUqkiqkX9IzbI4PomXePY866KWhARVq5AwAoIpPHj0ziRp5/1iAkXWcmbJ2h85gsO
wUEi0orQcAgL+iDYTBNkS65DNybTCA7UcbLx5xz+5ptmNOK7V8UFxCYKDlgxF9IhD1u7oDle5YHc
afvZKogKC8iMkTu/KnOAdOtl709wMCOZU7rzResdo8gkX154Y099NLE770hXT07RmXRu39OGEfvR
EqcMv2SPLRO0tKAoGMJmNiCVMHC83ARL7b97qSz8thcsIwaPD/mHfLksaW4AN1BLLS21tOxAKgFx
wMrPe3uwY7NwLy2w80+deIJ5TBXqa4O2pkup656OUU1erQSuiouyQGDdGKJbJ3qA0xNWwR7TB2Ix
dGi6U1fjuiD4DZb+FZCw4juuF/2hjVj/dtLeJEpn97AUtBteHod835Y6S1bEKVdeHjt1QM9LXgjT
BE1+sqSCCwmd6SKjmkZ/KjPoFnsOZEJnLa103J1k198MFNw9VnmHrnXdzvgFI0iIsCvuYDat9ghx
H5FnYR+ql3hK4oid/nmeghElKDgdKUDDlW/967+4TYhKMCAEcfJlP7mfDegeCTNBFn91KSMEpoAV
JfQc1bPPue9HirqIn6uvNgF+VtxJfU7M/a+ZkfpsUUlY6SkEgQgPIupetnftGhTHAdqvc/ccMqQz
5lwHRXI66iSb4DPrxDBuSxXuYaIHGQ78CI/nSXN52ieLNXIMuSoOFHyAvNc2tyDCd08CAw68BoUl
vviWsNEiVHcVjpIGBDGIkKM72JKKkk7XUayC6pORbB0Jz4mq3o8Y06kd7HID382jtIF7ToXktcPW
v0RpqQY/rQ6OLXDMYt9NE58RPYWfMmPtwjSXsAy74Gu/GVlzZ8d8M2oZCjXRUJS4Wqjc1X3tlqRF
yRj3EKqWHGuolubKdEU9SpAe49pRwERk4IeJEK6YTGfv/H32fq3a0PSHeV35YN40dGglwUI1vUKm
kUwagzUA4083XqzWCHC/jJBKaZ0maK0d1IP/IKbpP9LRegzN16jvz/bWk3FeI+aKgCnnE7+G5SFl
yZaV6uQA49/t3TiMV4vOaWYssCFviZOAqMs95yVT1Uw3G7UbQfvHpMbqoodn+YXmJvzJUG/ml58Z
E8wShR1S23JnE2u5a8cGFXiCa4UKN+B9043tsrKai57xTEuLS+kUFIdciP0p2MCZAI1cL0sPm1au
QK0VqU72jSRDmD7g/o0te1ttLDJJ01eEvUDN+vjAUFP/05m2VwuZzhSvQfL4TUbWfha7OPTdMnd8
ExUQjPvyDMz0HBHZU6MtTN0O91tdKYeKDZBiojPgMACdBA1oEcI0c0PYMwEtp8DmD4mswZghTF2T
noF4dlWNT3CWuWJ7M40PG29FyiEo5YTDFJfL+physmbAv4FfowjOGdedQxsXhngwy7ha96DMsTeL
dZQ64GESHNmSrvT5dI+0E9qVI2mN065O3wX6KoxNy2leiF46fgSgaItEaokYjN61UXmnvzccWZF3
rEGdPYp3pZEpUjg5vlMtvvzJ1UOxmdW6ZN75bLWWRJPdWd99BPIa76lJviF/+a+L4Z3XuU2yYEi0
Q3AIqv7Z5xpsuwNKOVqqdiciml/bWO8XkfXhhwmPK1wd0NcYugA2/CnEl/93SWoA8xJ/jQ0Gut+o
tX+hLVCHz0+LBioKs8UkSXYR+YjnNqQF+SqH2ESzKpZGf+3dJRKQlh3lLdVm72o9DcWfLUKulpTo
HjufxQNoLCTIcjDWPDD6VlFEE43M+BNWxuSXq8BzOfrul2IXyE4kNVvuoCJi0AXwcsiASgNw74nc
jOTVU09tUCG74J1Dwx6YSN6yz1TA0q9jiwnK8Uu6L+Qvpv/AJSrm8YQ+0VUziMWSdMjnKGR9bk00
t5nU+G8JqzNzpkS16Phei9MMoBai2XgKT+q8yCsg/cPJqQIB8EEOHc7iPCExuuh3lBKLLxDLoou6
Db1LQzAgUu30KCl5g1owZ/5CDmp75VkLGmPByHD0kBTz8Jdpb9YG+PWgwittwL0hK5eV5Aqu3/3T
No+8qlM027bYFEeO1NMG+MyK3FR16wjc0frz5/W9t/SmRibOWlfMSt3mNX+/AGynOTGQIVq5lGwf
pkH8sgl6zZKsSa9hCFsNbC1WtFiWWOogte6JcQsYoylgoLGdZGoQCTHI1KrVHlaWee6e5FZ+GLuO
XVgB/Jaf2sQmYtE7oiAut9FaSi4T+GVGc3ZoB8G5fOjoOttClJKKwexF+B2ZVdunt58NT7+XRK0E
5x7dNwOaS0PUDVFNzVstRY7k5AVPi5jaDZKiOlUO83DpXoCxWqdBUBgI/K9zoGHbRIWf25F+Vwdk
50QgjyRiIZsj15CKNLoHRJgwe1+F6we5N9dcYqM9k5xghQF8u0L7vnjO6p1QzZ9fqN45DO+WI0jN
j5f/gMCZhARLdjHNAHwAwacztbRar/j3cXMwNfW9nC97RoR2Wqd0PqqYNbte015UbYPtIEOjUtI1
X4S2mmYGtRqBfKM/DhvU7ALZJq5dw/jfb1qIWrVa2ZBYapDuBlVbfOxaHS79/aEoC7gre/agFJ+a
Wsxe7f7kNzaMDpUdcUI63IfmLEuWPebk+oM+nYw5Shf56jrIB51WbIt+OR05X73BjnGMFUWpXo5v
SI5aTDDigNH48vfmA8cyh+DUB44nwq11y3Hx2HhHi4qwO/Uu/ZRUQK58Xbc7r8wPApRB/QiFe0JZ
xnPqapn1tsAnte2SCceQtQrRLqz+uQ040a+MBQravJM0Ned/YdYpqmW0VGosRG4hQrnAJyY+f49W
/xLz/xhKhWijNikxn/nyewDYs7kkFmRuGsib25SR37R7SqdY9GyUWTEGSAEcR7UI9UvDyPQBVGsU
+ulxAEDI15qPOUt+15RwX5SmaubzqNyrTBS32jw0SkNuW0L1z+XuIosnj6/g3D60PoXp9Y6LFSCk
3kppuStAQsEIbezfd+YZHk0Cs+nGYBcXzqmxHBUDyx12hjRTLzedzfeET7LT9XJ24hbTAarSj5qo
EqS9kBO2CET0z6vWj+D2oo3cJLFnFeAKyhjgj+gLF4DFzhc5Mb92U/ECW/c6OaPXu3SdNpoCC8Ew
6ioqTOJl6tUKcieuriLlsnM15Rj3xYdNLXmqB6eNmYW3AEFczo7Ki9i7RWV4aZWzdh/p4nv31S4Q
DcrSYznWepP/s4gpSVfCUNnTToCRcy1/y3Mvog/x4u6kwVBHMgcHTAgf36tfvAQdN/8xJMXe5zs7
vFz6G4koYGdqPJdSH7k8eGBw/vuEhGCbKRnlbJTVciWutrWrdV4ZLw+dw/0oQVRKF5wzWwTIZtUG
8vaf85V0YMg34mGPhN1ATdWkqdkSWHev5jgoCJWQMO/4l49Syoc8fmzwM66eHPINcdA9hfXIaMvV
XXOoMKD/f7nF3CnVying4nP1soiG+FlCcYp/y8dRvpZIB6eH+17/fpGYt1THbXLnRuaq9EUpo2pv
H04cimr0YBjsM0xaF9Q/zPLZ+Cj1rQuBo6Z/lc+RIP2Ncook26UCi3W0y4wBqBezbuG4fKGIreUA
TwUw/gS5UAvPdeXoaMcKwiIRGj/zRJyrNEgebBWH3TIS6rkOWD33S5Is1s4ZOWqi49MhJZaPqlio
t6XUgPQ76ZhmnrEtboi1s4exXzCFDdJ1KHo8XhkZuJcQARKoTSFHchcjHQ5t4kj4v7XcGUJtrieY
bSAr064+u/QhZPDr6vfCKs55ATyzjjARpEbBTTeWUSgufziKDNjv2u3AdvTQ7k1CRCHYuf2veecf
oaSKnYcCwzT4SK1UXdML3pULrWxMR+kX6SmLLbqm+dsQeEtJnoI1Sum2LBdpMBgxBjNeZ+szRgbE
+FHrw3EIYAfleTFq0UEBVKIJ1mRFS81H+McXhcVH3V36LUy7PZpYivRH6v8IFQhJFq3gM0hEbzyP
NqVsxB1L0LUvO5illiI/yuGvmCJU6ny/uM6KLWkCkqWaGQvALMgrcdMrIAV6umGGdozsobR4abMw
tN/3q/+lts1KyLhBmbRvU4TRBt64i8NZWoI/J4dAev88JkhKmfwVgsRaYYrz/E4fI6oRQLJM7900
rbrakGJbSlfJGWRLiHJD5r9dRdxb3fplrhZ3d05RIkSMg8sYja2hlmF8Dctl0h9uimJ4MNGMPY3P
zVa6I7JiFJQB/p2Y3DXdoevvYq7VpDEKVGWAaqXKpg+AMALHMdp6CxrTM8oC7Ja957Y15GUtB6qw
k0hyQfgexJijOCgX8V0x4gfF9tfvD+BSmAGwqHIUqxSqqaWUiSoJ8hrQ/ah/mTunA9i2T0/I0/g7
5t0ba/d/X9I2ocmGqqNdgGdrhUsYvG1NdA/O6k2XsNrjtIm18p8L/8KMvOqvYBBcEPZ/JQxsDa85
6cXgBZqkcCMz6+QzMwjWKo/dlb4rjdZIRT2fZ36SfMaS8duUgjDaZQ9fNw4KlfiqLrjhH8ujv3/C
W+mo8XHgiW9zVRvLktUy0zt3eLcmHNitN9ERhTEkFPcpKRg01FeqmxmzsiEFu/ig5S6aPun37qQE
LR0CiBVpD5SOUh7/UenwOkONmCRko8QBCHluiGegw1KO7jycrCMomobiI6AGO1VwQnfckR+t6HvX
wprvnn/Gqax6t3KMFkK73nM/zk260qMgcb6pIJ2zLOWEV9A03b2w8IbW220AG2HjPnr48VFNh59u
G1h/AEWtiqlH88jYy00WyWdd2/moje/URNPe09gkJAuXSDswQO7ydLL3V+hMFoGERlgeUHzXMIck
oywRAUB+J2GwPA30rLmfb1RH9I0svry/TZIl23+eoCRscsn6uKNv9O4eE7LIKbVQb9xHvUQpzAXd
mp+XnHKa+xKJJYOAJTzM6izvzslQkjc/myy+QrY8GPF4Nf5Yl7vc58Ye+C4QIbuckhnYvIcvvbZ4
TIG7g+LqK4bjSxAr1Iav5DHP9ITvaSNl/j4NgOVWdJ0osOGdI6BpUGXHlxycCQM1zfKP1fdK6wM2
jUtSUQhiO6vJFVT22W+ugcJKN2IEt/31f2W3ZQRH62GpYu8J04MXZCtS9T9V/zSqyv4ekOnDNb7i
p3WcF4yxvgMlaWuYmXFF0m5bvJm/JsITfaZWYt+pMQ2sWueWboqqN0rmT/hofwiFVVnfYyQkOk/0
9IvbXjcGUsFnNwl7rxxCkBfZIRBN6bPpaP/HWdoFlqmB9XxYJuJ2P1lA1DyRuKN5+geEi0VVzKrJ
0sABu8ptFveC5+eQ9d47xm1WvQFgOSIpocWMnckfn+P/mXWdlJCRZ7xxA2LnXzgvzM9RG6AhEPpS
2Q/MfMxsx+gA8AAN+mICOug7UTwSpeI8NKK51T3tt8mTkzmQ71Yg6ipEvnK1tYCKmAdAYacmtQdx
+V0+/VthmgfsZlE1VFBYzZhirMGmHZwofSDWb7nvkg1jS0kFAgWb0MWgBusOarfvgD8l+YppnzXb
FsJTTe9xSivcoZgMa8n5LyLAvURR7KJi/VtGBtWbG3sTfOjWEQJ6sGxCI3qRT42dH+YkG6ir+JDy
c/VJPHs5ZkGJRyimGK5hdTOnwEhYJ/d03lq6wg2OnfT+nb4rALNwGqjPudBOT3VB5EDqfYJeiyrK
96j35xlvvRktg4lYoMfxavFP8IKp8mhmd0fizQZwWlt2tHyu7bh73zVFK1N3M7IC4WE2zTWpIMrJ
9rT7UxxKypYunLnDqb8/p/AggTJ6waD3ere/0wSEJp/Ln5Acgv+d06tFW32Y006lQbIWd9K96ABG
lOK2nDJ0xRgGSy3+GLSyq807AXFv3O7lp+yQP96Fn9Bd2IxV+80MjsRhfStzHAFD/L9UCCRjL+CT
gTUz1xBYINf2387tjrCeY948MmhM8K2igC4EGEuPQ9B/rkjqDyPu4W+HnalzKGuD+ZvZjgVYfGlW
fmKSm9jEfduU86q/LH3p51FNVizCj6VUXLHcbieRaRFKXPwRNmZHouQdrKdatTJO7MDbnDdvwo05
RvHZKXayko9gKackF74QjmexOTXWdJgWwCFFgDjJcKClKflS+p4hWlIj4jE1umaWV/xvRi6ru60D
epP62oS11M+Q7n191KYJoitzLLkGLLHAPHeevETJA7bWoYWPR9F0ccD+U8hBl2fPfQfW/1YV3Iw6
jfvQeviHvx21rTCKCPBwZppw96TCKOBhANqUbEfhfZCAGP4tFDxIGGxPJ/WmkLif0o4a28d+s+uR
nTUI7xY45boWqOQ721VTg04D5oJ55b3UT1ezJCwgEg6t2FnASkVkDDyGR34j2OjroijhCRnQk/ke
pddddXNnTZhdKYPsOb7k5T3CPFqvgtCa2+U/qnjjAsIVoLLDlQ9o/6wQBKwkyYxsMwN8ObHDRWV1
FbtuXjegZ/m238ecdAsZGlSHLycYLaaxhObj3+Lmq6wLngyvEFqe0Wdrmr//ttCWB+UIEdYpL/uS
TGsIkp1vx+WMcPvmkR/++2kEMss2dXKwvPUINS0vRf7q1BsG/XrSpWLHy320mCRyhkrgFuYTO5BQ
RPk3/qooijQpzUV2vucW6CxQK73dlkDbrO+8n+o+OkmTdd49ApJDwvqEJBn1c1RXR/Ms/Z0th2zV
Vdnc/FzTqeYLYTqE4uoCY8MUWgB6HV123TbvAmmRfH+T6FKbDlVt24T5+fCu6x3rTw/KuxV1Khw0
1nBk9nuEna6huBbfuakWwLy1oOfGrZ+2DtRRu/6CbebiCxEMPLW7Vecg8iKIsPLxFmN2Lwalkk04
Uoerv2GgD0pkVnT1veEU0NJQUvAkuwVS9D7YkNEfLoI6qh1hiaePUJWD5k1p6nRMjAYX2EjWpIny
C1Ol40ktmI1CT7J3lDQvRkNy6jLHnQYz9Ikt7TYBp0KVd2DWrd6A2Pfs/7Txi2BTYmFY2ktpZZEY
yo5IzbhJxYFIRYMExgmkwjWazlJmrma3aLEx/lSnysBK9xiPF9yj3Pdj0ktfVhyMjcGtjKVzfhFo
75aW+tfjvswHxT2Ab6EFwREeZaMLvScwymz12wXwSG46JojISiBS9mbqOaTcTnMoVN3ROIfROI0y
e5cqk3U3ouFCeC424R4+c2XUaybwP4+7ijIMuZh0sqbGIauD7zu6i7KGdpGYkCDJ4UA+URLF+2Cu
etHP6gclilM7hsY0OpPtriiJ8pj7P+0IZVbv6biUr3zE3Irf14lvnR0vd+EG3IWHH7ahlgsvPox2
QHKVxcQZhXh+m4zLmxo4l3SsE0Iw33oeyYn8rhZxCsrJQDPKsp68njgo8GIyNCBN6U027e9U3f55
XpD7uTS46Jgr35ylFqOkUGNpWXZFEOdilVHqk9yAca/9LO0oUjQDZY/B/g/2umX5p5H3R4HJUihq
BWMTrT6dUqOssP2vLHUMNjB9oEUmBj6yjRJyLh3ioohAU9zBZ7B4Jr8XUZRFDjs83XnCEve9htvT
Sz4TCCFN8lp1PpjR1Ym0oKFoGNkBz7JRZXlDj4HsJrx4h5s0kIRMtTWzMXuLYvqfYk5pCD85SrWA
0w636xqzkpy9KUNo2qy7LvfhAeh7D+MPeh170/a9zagGlZ5nLe+BTG1x1HFAqjXysYYu/X/JOIym
xVNY9DdmAeY57luVxpaHKP8QVajcPY4nhvKWRg8GAsaHhGLkv1pJ72xI/TVv+Wr0kc6NZC5tkYDY
8AFrVXU6tkCSk5x80JGiKiX+2wZgrxojUbyI6SOjrbnTOgv9A+W0/vyocCvly6wo+mxr2JjtaZJ0
80KMReEdPm5c09Saz7K1kWG+PoNC1/RqvdfsM2B4OmZ8+rxjphYi3sXGNbKZd3z8zAEWo8tPnKJM
WAK9gM24DiCXdwiVGKUuV03v0/F5b6O/Qp226L0H/5S5zz/s4p3gAbldzvSDJWpXVdtCaDdUGsqD
aYpIJhmPQtFqbL3zVgq5eQDc+rSlTnhTwT6M9uakdO/XFHYgqh6w4cmQH/CUnDUkvY8oBqHxEqyP
m9urKAk/muSGsPatp49ffRzCNmr9MW6WbXvqVKiKG8k6lMwfWgTZIJNll6GYwUo7nGWCMihdv2Xv
4Uv9bBQw2SFx9tj14UNmmBjPpN0k14JG8HqALuxc6AQoMjpkJQwmaidOs9f4Vq45Z6bE5eFjluuh
I5Lz6CMcTvuv9HMNqtvj2PSjrrq0h3LeQzpuP+/LHwyWK6pcE34JWWJ6+PvaPfCIZX45F27TyUAz
9zUXyc4vxFEIq2xTH0ZEK24TjYKESp2uYrtNtpwka6+aaZB0kwQnmWK8+GMF5jAPq7DxblNW/GXH
kSZRaoEhsgBlozi2KEqkzhZJ2KAJ9I+Nu6mw7q76cSZpGTY3GSvuwnICzFIcAlJPYB1ntiuQeRFU
n2qKM8cTYJNVycNlFVETo42AAVPoWOCs93YxS4aIesm5Beg29glXgJhzID8LVZzucHbSQn64F4ZJ
9Eaa0TPC6yTr2qG0VatAQnYBA6/vFnjHVQL7HKagSkjXFPVdzOIie0lSq5+3C+/9sXzxXhHJJp+A
lN79hxQ2oKkIXKm24wxIP/lc4BQac3WchzMJAUSI1EihvKTJCctZiY0s+7snNDMHEZoFp5Kw9fyb
WBP/gUz/Zc+7Hl0iUCR+cpVYlaVwHGsQedNHgUUocxMUky6Oo8HQ/PxGu9ohgko2LJ0SjoDGGu0O
lGXmRymBltsiTjocgOFCHSMIPHLwqhfEyqHJD4wgojY/hXdKN4sLOFkCWc3cYK5m0p6akiRew1EI
0oViWDikp0RwfeT6JnUhE9CHapg45rTQ34IQX4Lz4XVd6Ffjjw6RkI2oKIguaOhjPdEDq3Te4mMf
QjjIuq20jhbXAHZzqzB/OtDgD3I3+cHjLclddRlprhS73YnqLUuCUDi5Pwx5nyUpIZqwcLL1f1Tn
ZCngki2sgkDKDQ/Xyo076OFdXqPHd8DYP9/8Qw2jRTw2bYUuONzy09yGDLmNoHW9PVef5rghyoUG
z6lM8qTm50f13qfRdrfa6cywKa6jE/xNaj/vfbmdiKTZgdi1IGlZ+hcCPRmm5QnUCv88wxSn/W1U
iLNQbVLHMF+ACtYgtSKSCFlWMm1lqVJpaickY5wnLUrsei7QYekgaFiTXhcQKSHdy+VX+ZztiH/1
d9W4jMZh0cCKJ3IfhwaKB9r4h8e8DUMOGmH/KpC3/MjtRMlvqqXXZ8KNo7HzTbWFr0M1bDjjuWvp
IY9B92KJzxp+5f8gDwjVbNhHuDcl2wKwojY0CMFYui4QG0Y6ps4b+kAQeKqhiBGiKySXgiN+01af
iRsJW3CedoGlBSB65wEKvzMk7z7Vp30WDW4yH67eeBj4epaN6+GZAL9SrxNeOy25ADbLoqPurygD
TeLaS6CA7MUQlM6OYJSMBxSQfUR/SzxF/EDC0QGaoyQPqu03vVmxrG1xjWtORue+6tyUNSRcazGK
lRFuLfUKqOKFHlRK3y9e9KmkLm3MHDrcZl7UqMQ+zqgrfkpmrU5CymcHV85P4BCsjXwjOa9qJKDf
j9FI3thUJV027WX4zk364npBpFzBZJt2UFtZeL4sssJghN/J9vuie+FR3U2nmD6xJt6Xl8dMSopb
KU+/Nqcbr4iQpAC1LHP0NAFIqvArspVHiWfOQUuxkLeAQ6ND3JAHglCn2aQXKYLrVIl8MWUdLiiS
SvWiKcvr0N8t6LLjFBIQY8pTNlBpwydpPRL0cdGZPuRJEkpXlvGR0V08nol70VbdYpG+JbZa2ZLh
KH+ZooXRs63SLFIuQq7XoTclwCvAfaOaFD9HhOMNrakFFbGbTqk4tLf3nSuEOp2MXU3Cn6+JJFrq
5Kjpc4yTClj4QqAypSRKYq0LH59xMIB4yDZ6OAJRG9rCz1QWyGaV7SAbNORmFT8FaABvM8VOUhgR
bSl7GYFKhr12uuRh8eOJqRqXNMlxbX4mwv+VizEkRVlBp8wQQ9/4Rj+pN6fKAg/Xg+bz4UKnYJ98
x0V62TXFwQPxVw6ODw9EEo+xQozvdpf0sBp2xe+VBasWnY3VrAlbCDrEDDg9mzIpaStH0LKsFMJL
QpviHKDtqsa9hyetzUFLltiHm3nG+VPf/7JXZFbESoibBwVpanbBKgS2SD11ZQC7BYaTx3piBcrV
+wxznZZcz7xsMJOKLxZIj23Xb6EkplNsai6Dqt7TKIOM6yFz6DQHhhLPpFqVgrqFrbGZjT4pvLus
9DgmTFbOzYiET5o471Ued89x/kaanLoPpQe072o+tGT3IU0owmQDDJwg8WMaQmqUhXwLKiAHLXra
d6J1cXLYcRZmISbZWmH8awFT4x4KXRtjMdpfosLf2Op8qUn5gAk2S/fjLdBLtvlhIc5GzVuRbsix
k6kKvKV3HBOG43Bn55Nhy06dvRVfR5SRw4nrwM9df+pG7551chHYILMz0ziHFNFLc3F6mu/mbUfr
mJfS3uBs+qAj5/bG3YbeKI3uuV59W+hWhAhmfBih8nqd9NaGGz5JzF44PvGFAMB67/AjmMYugQwp
q5bY/v5QrvcnSn6s2UIFSPRO/Wq2X56ByF6H/Q48FV/U40cO3iX4loBR3EBOU9nmWB3SXv1EgKze
Zr23XvyY2vFvs/2e1goqlMtHMUyYVXqrKv/py4Nkq4Ls4zt+4OxI7XLMD5xccwOtt10xswJWC3E7
CDhvZCZyaLSBOfjfBSNkPKdPDL0aYnMCoSGNQwydfZTgL+fhgWriAXEiZOQGSfack6x8gjTJ2Nko
fEkGDQvvv8PzOJTXwOFCnjP46/z23LXR+1hAeiFepqTKQGBUMZRz2n3AaBQuvrBCSRl5S3gNbn8i
SlvjEVEnpVvvBOD4/1pSq2ctdvj8W5jc3MGQL2FILHhvT7qQvrjFvk/vtqGvuUy7QCOMk5F8wmFW
/ngNboFjiGkKPvRRlb9l5iFckr62rHkVW+rV0et+XF7q+8+nMql900K/SMZiC/7ROAN67TLLmiLD
sTA17JA7HcflsHF5wIO1C/sGqT97xOogeFVLK96w0jeWmcP2Bg+yg1n+YtelSrxkYDU9je0DrYFj
6o79OCi9OMgZaMo+q9igxitOAqodnZsfu+c9mtUuuO6v1czYqBJ3Knnzv4zQq1o4pn7pDWDw3SW4
sTnZ91X7g3Yy0VizuO83ia0m6HFTnrItB8fjVU+elAylt5e8+9lo6nvJRQdmfDJ5f6YTSFqpAF4l
Ar+TaP5H4d1b6ZWPOrjDze/6IMOSfFY3hHSDDjZFlmr2vIElwDH9/+6pwG9TeLpcgrGi0gHac1/+
AHu6+FtlCrW+mfc5gw9N6WAj7TzGhKg/GVOKv0+4Fo+YjWNEwHTaQdhyojx73Dtjwu+rx04kCY4z
DoQ5959WR169ipsVwyTLaUSDoeQmN3e1s2/UXtOgTAAasQYaz98oRjwyKgG+jcu3IHFsrCWEtdJu
DDewyD4goQ6LysbFn5kobXuJlItk+WENqzcSz9OR4SVCUPIsOE9S6kDxr1ve4v1stIjjmJ2qR42s
YtDGj90dfL1Bb2NsNKAd5M6L3py3pfMVs8jpIGQrw1jctNlnfoUKu+i377vCyX3JcaNFn8oVK8Yy
zWzsoqn4in4qMbVKIugnaVnsdtra2mcGE+EqrbUeY6onowbFR3cLrlMqy1yBKFU+5b9eCqC2e+7W
ldsaLdQScrsJqI1LbTLHk2Es5xPO7dJSOSiMoWmI4dzSHWB+pfWheLFrxaTNDesy9TWx1JH3Ymlk
K1/ferhzvBn6BrIE4zeSTnOFythIM+1f3jn4WQZvzknmxqGNUNMvlfl9nVLZDWiUfSBduSRQ5Gc2
Phwx9R5Ow2EVnRw8W1Wk6epuOxkPsGEV3+HRvcXc5kNzJdXSQQ/l/Y4VljW44FtbOo5FfDj1bUmm
stB5pmqX1CtGNjFBdMK8hmL97b6x7jayV/TKDUW9OXTrsggjiMuQesvBTfvqSTljn6YYAcdcuxiU
gUm+83ZoGFvc2r2rvxV4YNFdgwq7zjAeh0y13N3eooV2VYvGDX+8/ew0d4ytQc+dmNz7m4CabPyp
yrAB0cOnijsizeAV57HMOSB9zWcR1pH0p7fmK+qIQ/HEVt0Pq/1mZLHCO5/bue+ojugeQOf2Tixr
UCEKlEWK/erDqBp0eJCpBhO4jcdVgBCVhHHupHTVkcqK0t5GRQ8hRn4ZDRuU5wEBMjXmAsagx2r2
gKsHUkRroXCP+S5l+1WLuBMYFDVviXpYyCXwOkdHyt620knhxP/N/do2fsXUWP4jHHrk6GTpUvy+
zzj74XhwBt2enptpRiEHrx1oDJrU87wzKfaTaUEsdRg6ODXwBH9smImQnIBuBqFtAi5laVbIZhTg
Yrtr6/I7MEVui9uyzHLB3pkBEKlu7Bzj88Su/U7WznqVbOwm8MQlUQyMf9+vBPuGar+x0XW5MaV4
D1Pe50zm+29OUNm0aTC1fZ9VXyCVhcyTOrhiC3JfECrtQeTV/YzPXr8PqbLWwGbP6eBZOjOdoQIX
TxrGVTBVoYcvN9oRa2f2KZlcX3HYTWb6HCODHb+iTigjh3J7VEY81BGbtbIT1iNVVjhIj2fl/DiI
DppNuG6yQ393GNbAks0mOy+mqpZcldJEZMiRLYk1M0bSgwOpQ1FLwvzeWrt1izGCJbSitPPt/oNc
qkXBe83qKXWjqYBph4zDtVMh3sExF58l/QmJeKp0cYwIrJVGjaxNbASVNfhybM63OPEpWAI2b19D
TEUH5LUqxd20MfM6J4pXhXQnVnve29TQA/aQqglwajYBXsn4NyGILsscJVCl73tl/rO6Zv3VQHYg
udh7dQGV8KYVFVKsQ6MH+2ZQ0caapxnqpbifqCA90hbb0pn+dNcUvOpugrTwwzaBXFnosRRWA+8V
hL85Dv0u9LOAZ73T6PE+mJZBG4D01BDHskBAZ0Cel/JnrPLs+5qx8M3RKQ16IweN8cfQeW3lcMmM
r6+A+rrAjqyZIvCBovH4q4nPDabuHNlVRSPgww0AUpyWbcx3PwefkvSDX2/paQjUFZbbOiiyRuYQ
h9DcVGO7hDxbTWS33r276SphSrlKGsnAJQAjSK5k97ShAVuwoTh/rmzYzDb0hkNQFZDX68CNRqxI
nT3g7NnpREZ+EAjSffQkF1lLgLb7qTHIBlGP7LabuCEa2trcdLpLFpNZ1wN4AHi2KfXQtLFVHuB6
dNx4hTggis/KzK9KO/eHaLkNaMtiEeBj/+A7uAduzrZyISFdwe9cn98fsXURttj7lis2SRecfuWE
HOqKxaOuqFY2r8XMvEEySZdranimmuHKwtxllnJHN+w/54MuF4eDmZ7Q0+7cERkx/Zj5GWaKjZrX
U8dKUtaSMU14/c9h47YFdVvwTlUedmz/Vmck9YK1cEDTEg02P/Cpa66cx2U1x3xAwjE7WI40BF8O
YDyfL4raK4mqaAV3ESGepk7qtVfUTiWnZXUVJlACzouegD7WOU5fwDG42hZfcGuiXzX2k/n8Abrz
ZZ0vecPLL+fuR2aqAQ345LjOVvOsxUIxZwOVEsYQyE5vG5/lmp3ksgpiwrFhAdJJ4dTL4QCj6iam
wCZcPYneD+D6MfZMepO1wGblt4PTsC+yyJHSZdbSu16nNX06xQXGv763T+Tuso+oViXu8sQBYnUj
ZkICgqJMh6stxLYEN5De2BYCdaYCkh9HvmrO0We29OgbRGd9Qv9JVHUnVs+i4MscYEHBcMrFNV51
z001SHdvzU7A0LoSu0392exYCc+b5f9luCU0pn6foIRIJLfM2Ep4rtYDJI2TNwZLeU71h+3Y67R3
ckAzGdQ7g3NakomXxRMGqFqlpmB0nP+DGF1YxrGcD4ZfoO4/ClY7BQL3uYWAJg8QjgpZ47/sNjWc
xma9TStbV3a/7PtwWULYOcHoXsKyvZlp9FefUvTaGhWNcqjfTRg046xg5sNpp5cH7wF+b8PtLiOo
KfxdIJ+RRwdw0SbsSJCzDgItOowyxAX5hyMwQo516VmtD4gCst4cnYuSWjczR8GXYhAkN9gosieG
R/ZnYl8YysIDl0vpf46HUzbLvhnEqeQmffO6t3GLdyhEnfPGPXrXX0tRVTaeXfQ3RLTep7eUPMc9
g6FhuWvCcxPqLXU2vIdrvBfFBrdzlyEiOIvH71jQFpekiQgknSng7dsCpQk1NgKSdt5IpBERP+g3
sySVIRJIbkxtWUD04vNk567WjTqZ6PTlxD6TYckFx+Rvkeebp60GJ2xZ2BbHkkp9YBfHvooHGVRr
M4MV291Zycs3GDYuDxalLdg8kmPwAyfJAfwc49EwEz2noAlIRadlwK0WHiI2CXWK+Yck+tyE6B+x
dYxPxeEtan4xjiHi0TgQ/EPsqda/320mDk4OK1/YnUsxRO3O0Too39lfy//EBzy2nCSy2EXhe5n/
3pTyXKZSEvlKsx0eDkaaPs0SetJI2uyYMflfNVgW9MGHkojs0hOEhvJgEU7K4ztSaLYz7EjMn75v
NyG5JQ3r48vWuETMLzO9LEmkHHFhSRkG4Px+JZMC8bupjBveT13E/hWldysMr2fp2MR9V/gFGY6d
Dzp0nvKkS/C/vPhYMbayd1DqNEPwQbgrscHHtIK7MyIcRkksq+8qOuqWlEVJkr93ipvy/h2MJcph
uh4wmPBbZjAhVom3/yhIIPFuPEU5Tk4vsoTXIwh6zUksC8U/7MBAwoJedyKaSBt4nyFxVTHVmEDi
ubG0XIFo3F4ajrEbnbyHrECb8aZaHEva+8kkFyTJLTnC5m1ly3I9bnedEOfP7oHQaQTIO8858jbq
5KMUlObJ1oYR1SHEdd2HWYzjPdpmWyzt/KTy08ujjcVZ5wMRz24kyQCQdwvPU+TA36v4f8vfSH/p
PMgqoTV/G/lqZw0494SGAoDaG2n3l/EiaaNXOITPijzpWNsdw6pv4rXBdscCDng2PwPjnYSEbsiP
ELN36xPotNaKwVRtkGh7w/CemeZTPvgEAbICrZYgGX3f6bnX0FjPAYrMgSwdQdSa/+bNe/Y4KOYL
WzsKbdjh65H6SFgx/AYdv9ZVMjFFpQMjewXWB8sbu6uD5QukDU1K2voB0XlopwPgobljuHgMPGau
AfOfGzA5iJsNRCPInPLp2uZ4NTERgyTsSyxSBTHGWDDzCgegbCFEBzfHV1lwB90SM3t2nzMIsOyZ
63O/yrHZC+Ja+L1y1Rheo+jTHDc7qz2cXAgX0gM2RlPPfVWNA9dRyPc21H0NhR5qCYDZpribajFM
gkRP8d1PTwtW6tEZ9kB6diEGbzjFxxRXwMY5KpCVjWrieHfXWdT0zezKPwMpY6umeDx9upaRkkvn
Qe8lyD4eQwvtaM3CFHU4MfwtZnJh+p37Ouqe4Kmg0bn121RBTXHKmssmKmJ2zg/slAOeBM0TrwIS
Emn+GWs3/JWnXptg8W7/jY2z403XlqHh6yMOkJ/+fYEIxUILUdHViQd6MopnGn0GN3L0Ts8nnVxG
DiTC4clSpMHDI738kcTylxt5Afuf+isZPZfhZQ9Q2NcYxxi+5WOzUgdOnonAptIirYTNsKyNJLfu
VLBUjW+rULm9ySILSlZZxtx2XWkRBi8LuLB/u4aVZuuARjQV4vIwoEym8LHrxFrNy0aUUL9s43VJ
8yTfWEKhlXrDPPC1mqy/oo5xm4r8ba9Wiwuo92w70rA2WigZwNGeMPP/V4ay5D40qXNPgD6y5ZTZ
7eD5Comf1TRbFWxsE+wfYeINhNpRy+Nfw39qlmeOzoxvL4niY6NdTF0v4h8nO5dhrkLuWHXRIQZO
x+aTzu24X8Bk9FISFCTsx8sofQYurMF4BXbmMY/cgJasFjNKXkvtUF28OodahB8fvqswMJUOKYmm
6HHTxCZXKtFlfwbvJEkhQliE4ucFYku/OnnHrfbXhBfEpL2hOAjMoOyrEbrcUN4HkpVxyDFJTxVT
a5y+ABRS0XakPeTb2j5tRVkTjBk9guGwB0pvMD/8n0tlC78D4CZIBMtnm+/GBZlLyCfkUw/gnUAh
x8EpUV48gzO+wr6/n1hg8o+b/O4XQSWagFSX3+eoxaday6krfmF18wzIiR8ozBB7JBs8TosebzBj
A1YzKAbEfVaNjNrh27Ou2KSLR2z3uzGrQAtfTwY8GidSxJIg+1KIGXcMz4nBDR/Ori4jYdUIpjJB
t23APJlmOqJbkAJ2ovecEJoHaGgYiMK4mMl0TNjcs4mHc1gDZ07iD7TBUo+ENeh86KNyBK9Zlc+J
Ii1Os8TIe5JqM6pIqKpl5ElACnT2jJ03EbLNBqPMqUMLwrd41FERmNnRYPWA4qLtSQ5qfgdsIrSb
H/ucDnRpyjYWOiVAUysTc+BX75GgmNLFONnVmqaSbn+q9a0PcHYFJ6QRVYmSU6pe3mYXJMq7R7wM
FgwZpbMg7mCvlZ2qkkDeUq2jvnq8NiWHj+viMAagJmIkFyC+/n0+HhdORw7v60CfeXIL9Rqthvur
dYUPJ4U1BOmNAVxlN01MRqtCzyjgFvjGX8SbXFE7CrcUaCxt5GgrPNgRj9EsL6r7Muneid0fOYH1
50u65hAaYaFKiQoK1lSf+NZKC5CGHkQJmmDNu6Lu756TPcQ54eKw8hUcFt5UPK/TAS52/cmLELJC
uGCjO01i5YNLCfYAVvNN3F1acRoDpXNFxeOaXnH65cnhEOKTzzPG6dkoZp8f9Jxl3j6zrYOZU5UZ
7FwZfWoobqHjreSy9ugM4vS2D8BK6v2hZNAJ7LiDQ7VRs0A6IJ8c0/i1x9sRyzDu1n6xHFWD/K7X
jzS7O4A7Lencs8pocIq/653UDtGBvZJ7r2cl1CLSzNuJR7a8yfOEYNgSB/4hx683O0fEZ2CZSWL4
hinUgDaMG24FPQnuOPHuALgCZ3/jPhHmqE7Jh2mfYVpzdc7f8fo8wT/KY3cP+qHpdVRGSWch7OzL
5a2sOw6Xl0JHUwjWhqiaDJVXaQ01gG7NFVsY2YwIHWvIJnHybMLDcnXAzhcoueKRcA7jwyYD/XYW
FAT5tuJtPgIdjDTp+rLMZAo/PITn06Bi0g64jR5+19FjY8BiSE6eDiTPbHX6JxpSUzSIwt57gw5r
DlAcjNNiivIOT05oUk7CbtHeW+UjqFVHR7sU1BvIR2nw+RlPdDOqPDeaRLMNoh/XBnliOS3Mh+QV
ycE6V1X0UoRec5lHaTIrcmTdquhvGY2gdHV33iZLFp2rutl31vDRJpqHYtAr8LzJj+GBAKoC40+D
7kARKoMh9G5h9VgZjjqugtcIiQ+FmjBHA/R0WfGdmnc7snSHVhE3me4kuJvblb3q9xTd2w158KCq
Ie9poiU/TNWQRTpIJkrkmamARO3t5kQV8pgEs4YFtz3GErPWw7VRucdtkCXF0LCqFdJXrfk/dNIh
n3NIeNbbt0+YPwbIHUoNVUy5QloQrlWmgOrTfdTtmk9qrnomCOZs/QJesClDeMX+mebyidNIR+JP
aMDMMdt4fN/g2uUq+1YMjFLl1jHdaABNo1oqqvURc+CSuNrnmrbEAPuDAnza15ufZktYsqxDUpwj
hTmfn0R5NKW9TfVLEQE58fZFu9w3bGvuUufV5XTerktsMzeyZZhm47i/UWdGr1i6qaOGGrZICgO9
MJRjbn7WHTbN1uVxC/lmW5ilK7G4u+C9KaRc18Lu7aSV/VlxjF5JBdhlX643v9p24krPNN9YX64A
OeQXbttx+yRdjRVw4ai+TSLu9AIp9LHqJJskFaLRiyPWMpixmWj5Qx22Hsc6trEgZ+Y+rk6Jt4c7
W2U/tmYtrVNVmVvXQNmcCApLDpdsr8ei0rmNt66nugax9GUNY0UuY3mUxS6iHlffRviCKteQoivD
ADnQ/leJBrlpDrmhvybe8LUNF/EMS6fcTGtp7dFndaGdFOhODMEK36zvuxSOkT9UTTzKuxUQX94Z
k0oZ3RhzpJ+7clg0lAZgPBxvsqO15o2UP+8iSZCM2DsskK2Hth39qA2sDsA/38y0t94mxiCNe+BN
9rS09yKzLj6STkKfjsiIrVHC9pE144taCw76A0iwFmlTpPLh01ugDrheH91tBmU/gWNW27bQrv+/
cNXxPCeX8qpbk04ii4GYcwwTdLd2BPzq76y36+XU1YVPKrWfDSwZ9gLaZJO7J3tFBJQtUn/FRO6h
ed/M4X+hvkGjbHvU2KKAWdypn8yIhQLbj0MhKxkJZA3DO9UioeuorQ8OGSbB6bO/f5blOa5nNIEn
jHSI0A4gJtvo//SoLCbK+XhqEkYvaW16jPcT53Vq1iNuIn0A46Y8VbhBhnLjUTo8ibvhmX7o3Yq/
QRKWNhGynC+MW8GxYn/euKNaBFW11dVbmFckPMaID0xC41iDpEiK/+g/siQ6nSRq6UtIbmXQbYuf
G5U8azjhSFwkj0+N07TVm6x9zSIUveAhjhBAWsNfPxUV2WWOsq0Li92gOVgLOZ9w1gSOVXdi7aUA
pDRR/0uREa15Cntgsr2zHZbZEvXt4UhSv+PO1PTfT9ljCAN3uzlcRdBpeWNZil2lPWCPLKqXK8jQ
V8dNVLu8IF8BmixxIYEsYKEDkjNy1VARpiHdVsU5DMEzAOYfgtJXY/kPgVnC1As+WZYs8V8egeNZ
sJTkE/pi3MiLiZCfqSbOSoLEcXLsLuE2SMLNgw175UZIWcwxtzIgtcwDCIW0fT8SgYY7WHTPFaA4
erIlbPRCYCwjDEt+a/sm057AWW95nj8T/1/vrsybLfiPE9OJuGBcUBz1PGIbHVOnr9a63hFxCrzD
X3mV2vHyI4rnk8HpGk1LHYxoSB1itp8khnghwOAFqiWhh4dE5UEctPZ+E4kzbK0xTcGw4inSpaMz
m3FZPvpfkK64ttIu2mxQpxw0ZBCJHoC5AMeZ/w4vUvASf+VvmD7DcDcWqSKDLSRyLWwzo9q0HWPK
Oz1/cXUopUEDQhwyrjj2IEUtEvDBLcfq9MA/OMx3tZxw0Yvq5qtH5x/i1z+p/dsfojgrBR1AfEZi
ALBS2CC22PzoD5Jqj/tsbe587VwLtgnai87QEzqweEZ4C9A1NV8vb+R+d8DjlyRKHmx7XCuPKMIS
bs69j/xE3rXfuAhdEqFMnbkqse91gjerunQQVSm2B/AgiOUDwGcBEgg48aHuJKUAbkzaCwOXxXCB
lf3m7X67rtItvvFMxYUQC9xu+/X2NYZb+sXw6Xlvev2TI6cFp9emFimxARxpSVXEppidCvRJD/xU
zdQMfCyu5MZYtzfS9w8mEASOUPbsT0cKVuu759NzEaf2WlAOcOnQkenejSGdYNCx+sd0CUcWw7V3
SLVw8trnDLDy5DycruVg2eAnUiYqDb51YphxUtrz1xbjHGSqK3Trf1h+6q+AV5eWAgmAVA/Rfw93
8syACP6ktUDxZWqcLDtakphfd0Q2JjfO5KfQ5YQmk1maOazSoeM9FlgmIHgGEmBqre9CuXo2zowF
UF6e0bYtSJRT0UcgodP+BRF+TxBgQadOgC2exy0u3THCP8VT9ZFxbGEgtIrofrHShm9IpGgLGeJV
ULqe0/aKpr3nDIWI9j22oZ/gbnoUV3SpCyqC0+8/atNRVC3q8NQJiNvUHlWG0xEXycRMwFe5+eoi
lOloZXLw1kqqFPyHtHKNhdv2Bd7h3vGb31JJqMHusL6XXHS55FzFM7a/hmSu8tga2UwkC8f0+Lct
duRiOkoWAY6X+lOEgwm/NuYcUYA/mGKB1SkbbVHGnk4sxtnx4qrX7RyYjOssfqqrHpbX4l7brZuW
IX2QHiiRye0V+soSzOrQfSNbAO+wpfWebBCe2+9cAGUrgWzMfafYAVALDxLd4Ax78iRtpPD0y5T8
M5GjfwHbxhRw2GB8X020BpZ2BbpRuTspkl81yoOs7uIOz/4qKsG4EYgFeYQ1mauXF3+lbfi9wuDa
tzYiLV1Z7agkmTkf+ueNC7gCcowLSkPfSl5mDXuVCpE0VTT60BSkGtD2HW34c01Ygs9vGSTyXQve
cF2evy+n6JW4Gfpid02SHS2ffG4yWHTgvzPmr3Rs8R2lIYnb20yLHeFgYO//CNFxKCvMvfkYTaYE
rPoKGYD2o8Y6Utb1lPEQHS6cVql4tMMZnFNe6b6NkMLzx6UaNJNUYVa27eBamuqqTxKR+uNl7vpe
7HAchUBQyh4fFJJ4ojhkvSI6efgYfApIeXj0hwgikNKLDM461xb7yrGUFsNFcE9vawy1rRqcLHcZ
kur0fqerJzD86Rk8lGjrTLJcezWkmxv3pKKa0oDjdP7gCuwdd06+AniZaCyfbLNghwB+/sbdGgpY
OoTcaQgfNewx+ygk47zLhzI3WaAL8CVkIwtdvsZViKeHx5lzyFMPkx58z3W0H5D3zhbiZDBCe9P7
Ilmy7QYkubM9PgMbWLP4Ue9uZinjAukEky2z9FsGnW00WTdjLg2JhV4SDeiJs8mLV5Qg19mls2IE
A6JugZ0ppI3j4qFCndHxkRsjkpBuFUwQ4eNoQ+SlQl05eCPCWH+8e7C2EmUJ6OUjkQ+7BdtcZypF
eTrvSBGk3B44Vci7BtbmN+FvExU/C8jKnDnMVCDFmW6yf95jjmRGqoDBqK31ELp9A0sCdbuzn7aH
FzAYjjCkpKaX6gTH27dmHKxCC0dfpfUZIshqgd7+eWGTxMPHPuqoNyko0LP1WUhPzoyAmn+KLt+k
pdArYyTgyNCstTUkAboZFMnOmnlvzU2Zw1CJ9r6Z0MFRloQQ0EmB0KVDIXdnLEQD492qKO+NK7Wv
yE7PMGBU4ueF8T6p4Ba2tx1WczAVhqtLOVNt5tFVqXPweeZYBvyGTPKmsF3yMbZUqLACrdPzLm9x
T+0hqVBjhcpGJ4E3uhek5QJVj7jK47yvyy1ppKQ5tPY0Lx2GdS1/yd+Ava+K0IU86SLlihoneDzM
vcVSTwe1ccfm12vu+n6kA2KNnXtEY58eYlqyoSHoBweyETJqIDCmt+xCvear15QywNbo+Z4g6ETI
+7UJEFJKq5sJnbZVRTdV5PQx3NFn94IOKtRxGspRFpL8CAS7sdqRqOzKuvRQQLutOHhVn6IvuqnU
m/HpnEatyqEBeLMkI+x1Gag7Cca8AW1eW0sb0K9jSfFotZVDnNYnb6w/tY/EVE3QDAZIeTnKegpJ
gwl3o2P0KPotA+q3yEx8BFF6uGYCUaqWPMg6Y3vONP8D7zGZkufEdmqfM+IAhMdyoxZHjTGKDaW3
Pu6sq8u880/JIfrlIvAdYp9ZqXmxMnJRzuJbAp+vstSTVSp/Fgsjvnk7RnNEaLFyjgK1paxarEtM
2T9KXmRYOrDC9y5ErEUtGA+cQhUdn1qdXv60VgHAZy89QkdwaWYOWeYEP0/jFt1oEmBQJDbonx7b
7r1849rP2+QkH5Ii+WAgzIxwjkw15W1gz5xQ1bdF8fhVLo5yBy9UjSOL0Gmfg5qOOMSoKVjIxhLi
8rwKXBkkpu2daqHjtM4PMW2jFir1ijJ80+XOQXkl0YXPrAbTrjYceak+bFUWkkpLvCRToPiO0jgr
KrD1O8rutTpialonzWblCej2VHU4drg2vT/xmXLOaeJVLKZ52TqLZUCaAr176kz8IrYURlSx/n8X
JtFZ59IqLkoL6vyONtcfr6/zK5kZyjizP3rKBBK+lPzM1NKaFwzWn/mUCeqt/aPUYji9EOAdFKT0
gG434vAVaifcqnY+UCIcH2XwbukxZLQyL+WBrn+mhDY/yVkccV9znfcpcMUjZBEBPWEjfcZS8/0E
g+/b8LFwQu5VmHKGIrAyI59uys02VNwJ0wUoCX4vpI1A9SjAwkkUz/gzQr3UiBB6P8RfF+KjC0fB
FJ521D9nFTGJWggzZAHao4ZJzqFFUXorpyqoLMHoIUm2GJSJNK/K6cV5HLEHMJbaUwOGrZXUG2fy
TmNnfo0r9MFHQVgIspQzGKQPWuhk3WTKH6fgXbVLQEXsGQE+EdzanQxeANH59XWZ2TePYaWTXls1
22MCT6xdK/cCK1FiyYrk51qDpsDE9yaY7c4ScNta34/vtwaNhriD64NffLc7tV4V3MO5U4Vyu/zN
0cWSNq+2LFPCEKFpDcxbKMk0fBrFdFt6GX+MKrMxKfwS7ldXCBtQ+HWrMpAp9KhpR1s+kQX9fcSN
cJIce4NXn/euQ6mTcj68rglhMmCWflPd2irSEwBMA++GBdN+VKF4+dS148tSry7r8mkLTHYomrGr
E9092tLsuVRFCcdKAX+d4f1g8qMTJPEQwtZIpUZPihW/Q4AGGPmswqAwDZ8Oy5Q2A4alpr590wiM
DPBl9zAccebHymxYI9W3Y/uS9X+2r8EMvNohHtQeiFz3agidriZrUmE58FStqL8Qx0pRthBpvdBb
1sW9VVBAEwLd6qk6IIgN/pO1gBUdRZh8I2jsrbVFKrpGwve0uVRZ3Z263jCu9lTA5v7FdUVZJiFB
1vFiHXowZK6VRIw6ltifzT0ZZ3pL3eLfKs/kQ84WeRiVz9JXFMBRcEkBlvGzz+SF3/yqsNQQrES3
3pnOWGYhb1JJbZZzRwA/d+LvfszWMDt0dUSlfOhH88Kdoc+Od0XkbrL5jgGo0R8fcOG8mg5ci7uH
+xctOU8QHFD6/Pxcrpd5MBaKox4Fxs0FGqc81cIjb75fCTqPjOh67IjUTbHfARm2/Yhk0U42mr5f
dezPhyu+6qbWWjitkHgP5lcIWE2nyJVMpBpt48Wgs9yXzu2pdGLeSGgv9yLzy/VTmphYnEH+wG5V
X804GC1Zvp3prq1zfv2IllsJRgNxr+a/J8fkWe6dZt0JHtpQAg856gj8sXBySO2TXz2xCjlvOkVo
Ca9Xb9t9w3Ss7jgnw0Ku2ubqjEKrmM3ygISjLygIcXHKKhvXDC8qZPQ+C5uscENk/uIMppaEVGjS
1IDp7wHWxG9s38aniRzKeT0E6Ar6w+vX8p9HQNC7nWtW5tNovpoB1vt0S9ueOcabsR4Wp5fp9e0U
CKskYXroo+ynzs0ItHx6Sek8cveUOctaM6Erq8JL1Z4mC7jT8YdJRpvaC/byKYNi3dwfAczWiTBD
dZMe6EBJC+D+bkgAav9dqmDPA/Ow2YLYPLwDXNitt7/DGCmoU0YmC+5DEQDWC0qwH6RtKR067nFS
ltuSHCOQaGSawnz/d1SZOk73BkameMKu6EEChLF9ZVIPAaBZ41g2ynsFKI2FxJVcshw0TdK1lOrb
wynZ8CApvKFcY5r5uWKn11cvthndvCakornIJPPCAgTFCAN3PcQhzFF4zY/n/vrhZ6uE/Ars/Oor
UAgrr7Oe/VGHVvhsrAumwjUi9ysYIqgpK8lDRRRZIy+NoyFNji4CLWouXrTC2pv5asnRw1tM8ETC
97N1Q7ZsOkp2R39hOeduZBVWyKpTjNXnfqo8iuwIMhODGJjCx6cOx0Clz33lo9vrxLCtee8rUjDB
vD9P5YkO+2n+QeHLlwHjQqk1VBo+G/jaFsSSqKIMIJ5KQ9zrCoan5CNupyuf9DbisPouKPINu2Jb
5gE6JWnOlYllDwbKEYKnH9VAgVn9aUqvxv7pTQ/Bs/6d9cup93gBbNUg834USD28Mn/INeXzBvff
wJVzksZnNzJtD4eO8tcoHpLy/bQov65SbyAGu5rR1k+ET+FS7k4p1KJDiACmXaKLYvcUW/LE0X+b
NHFB+vfYCzz6O2Ffm/sOgxYSY9auqlcmQIO/Hd0ASfrFoa3916fA1MSEtBgfNPPQr/0XAMqx78EV
k297b13WBhbEzVxGTRFnyn8c25mVvcp2qhulyUsZp3UxKqqCbg1okZ0Xa1j16sJHeiigHQcnATvp
zjXMtiMQPRQPn4kVBYEZVoNSapYRhDukOYwgeGUpXa45AKGadWTtevbE1hi//U0M8NlcuXLlTam0
7vM1QEIMgrLMVNIZpHEeuLEAHkOxPrt4ZXLHJlwhvXgdttU418zuE6Bvpxb7UXp9JPLCHfWIf8PS
ZUZAssW+asO/Es03wVeQG3a927FQugz+TC62fztIYF8vhVolLKWSF1Rnx6et5QJkgu8RplM1Z/yo
htqq4MbUj2SxSdBxPOoeZy7PZT+ptEHmMUraGHDOZW2/BRmgjhm33esvFAq2hI0UwAIkUZ9VadqB
X3iwFgbyQnbgupRJQ62W7sD8EvB+h7daUDWWPeKAS2ft8cJIqjlCAFIUVBXdIWiJVYHmSaqh6OOC
EPNgBa7n589J5U04EmN8hRpXpzUowIxHajl2BXrhzgEnKywCafCnD8QBGSbfmufOnFjDLmoGF3RN
LorrZ6AOuVHGLv+jekMKXrXxJBF6KAyyfCY08H+TZ4uFq6Z89TtYKpZK58DixQqJQJFTgy8yZ8Sj
WADO0y9LbVxHtDWaysIaL6E7p1TgACJKsMNMhb4z/lBa+XdvEHDfUQXi/aO5KX2vSO9cK5bKdZPc
KVfbIip+P0u+BlFdeL9s/E4T7btWhmQyJsPN4bOoXYW9IkqAjIshv+jP0hMEFRFu1Pm8o9XblaYo
+zIDpjatgKE2T/dqGisqvwPL+DmPe/vZ/wxA8N7PM9xxUeCQertkjxxtidCh/3MhbpcW9ymtNGVF
zyyFw/9DWzP0w5XLsTgjmV5wNHnKKE/L5qH/u9fU26/5nkzyc50rTRAJT8J1eg4IfoL/Yrxeb8+4
ZSn2UuoDtz/QL7IePugnmoi00LaFqHiLDoxyjDbu7t4PWJa0Bq0irpfkDniTm6IPs85Ng+klP+CT
0j181tefnIWDHPaWz40S0DlL5qXIMANIMVT822IIPw/OSL/pvu5i1PzkDD4hwrubOKSR765wP8bT
JQK/KJhHvanCNRRGEJMQg5pGNMpUCi7dOTRrHRNum/WTgi0HUu35eHYg8a7Afn3rbLiYTkQ4mgRp
Y2LJs+LPyBwn3/4q8jrUBQCY3EWdxuisXvSG887lQfIaaQYBdjV8A3MF9hek3JUwjaRLjyOkEhGv
I8EyORkBaqbOB/WO3/F7hj7zCxX68CKp09TlLqe9sBwuVg3L2EsYhxUVzI0gscWQcGU2gywysp+g
cahvKGE/+D1WgQcmz5NMp99U5GXljquYMOl0rI3FBl4ZQH5I5JuSXynNAjEUXs6vzpqaUXzl41Kx
hFlCpVeIEZ8NX3s1MzOVO+yU4RTP7VVWZvb7eDh9X/ijSvcomYQaQk8zRFIfsuJfG3ZTuv+DD04w
cfoJFegVroTZ0vcLAFZwW1pmUFtMTScrwrY42U1fGFsf5HniddjkCJZkhYRfX5cGUEtWDhIes7XW
pIepy+euOoIbUasY3Se9/lyS38RdCab6JA+lP7CPIOPhxVta49jqnJwexqn9uNc4aLC7uVWJgBKn
gf4di8lqUGSaMy6tFSBX0v065QhTZmb8pTffD33HkCrK1Z0eXAiKA0ET5TN5y84LFvpQX256VrPd
80NVf0TmXtYz5O+8Il7Yji5I2I0b67WAG7asg5tew7R4LK1q5Y+VUdJ7jgk7z/vars7MntAxpw/b
bqLh9ZwQ7hMIgF289mzxn2h9w30ngw8Vls4kr0P1efQy3NK+3FsVz/J7ahlDTZXUaNBjyZhVl1xL
SnIEg0xzIxKsJN+HzHSW53FJi6SozsuFwDMoqpssUGcanxrwhw01TNeWpCXMhIXmejeUVqbB6jna
wtSIGeGS6c2F+v9yKlLnDCenN7JrHJgps+hg4+9HRnD0TDkz1ta2B3YYFhbu2yiBEyJEDwdzyzGP
2wKeXrFA13uHwJtXfT9RxneXm+O+ajOKWoYVQoQTAH2RFlKRXI2suLn4g1PudhcfHjOvri3OpwZB
PNc2P5WOOe8JsXFvVNWY8tMcRmWCQfwHhxL+sHqavHUh5Y6dJaCHjtLE1VJ8tDol6QS8OgllAR/t
2Nk5XAyy4YsgkKUaDi9Hp2duj0JdVMD9f9K/cb7AQ4JcLK40povnL1uS9cP4gg7PESmN6DvxysfH
xAAS/IBJ6seDMmf8q7wBgQGQlwzidr/XMsXLNPhpm0Z9yv6SAePctV6pQucuSWTZ5072qliXoavb
arUxjw/Dr0yyn/25DuBABR2gJQeJS7bTV3dEJa9JiflOosjBv7dQAnOU1PUuLEJQVNCV1LTo2IoG
vMPiyVA2/aiBXUXiinbRsvTgKSxXdwp+2HLCoWsfMfWrB5FZKRKWTa/dHast1oD1F/3fxGaxTTGp
5Qf09R0L6NWdXqFBDq8sSVfLxwAp+b7vquC1AsMhFUcN+XnSGnhOLC/ukHsh9EuOkvAMZUub5OfO
VhIHaCE9UKCsyW/Wl8u3mnZHIlN4ZNvxg3saM1g3KRCXMO+6pKkKS+dSEdH3rKyZRN5h1niKwGgp
PzZKBxpYgCaX0ykyV6cGeF58cb9HsVqVe7ly62y1eBL7rZSswbroNt20QcDhsdUbC2pAxN1Cc1QA
iSKucSMqZiHC1bYCQuke4+ONQmNhb4Ezf4hLe4fyXR6s26U1hZSIOBHrECqu1nTIa4dSe9W7XQgM
7qHGyaULt8ZrRM9wBdOKDEfElNpE2mUqBZ4Kuq+86YPf/8EOGA5RKYFkjnBPgPljYkG+UylNHYeL
jJ8lqH5/BDQ12O+gJ9JB+VDK9wxR2oxQpfxa00EKYcFm5gPDXrhLBOyBz/ZQrg1sQkANjRrTAtgS
0fzGqfd5M7pRcA1dtPGEDk2KOLQEaHYXM+GEMzWAweiCW4ca5FZ5nkTQptXkx3wl2P5STWYCHHPN
lYrTEwyu2JR+gxBYnMVEoIRqiK0ZuGGWPCRqePEmEcFonQzYziHGNcbXmcYH2tCLTfZMlviEbvGc
kq9+HIJwq3EtIIA2j3vAqSoKzgdM3tqKLCRve+GUJpfGOdDSpG3/Ll6omY0+ixdm0eml0bYZqawQ
lr1wMGP5RjxKlsGCwF6TIH7ax2msB07IBw+WbzdmDfuuKcRbZdFyBXYVxMr1vj9LzpR6vC5Kbja3
vN13t/TWuDMjxxEuz1AsvGv9M/TF3CPB0fStnm3Cq57BAu9EmHcdhdEkl7cQVevp1z8yQ3U879jx
sNnL6AJIrvGDwXZQRJDVnuuxJPWf1P1Wk4MOEW8gaz1bsqFNOIojvqapuQ8/xJ9n/qDihFPRCaIM
OSKetZrarv9zawP7y+Os81u+gluufW/h9Z6jYvEGcSdu4Uutg6Y4dMFAiRExJoJxHn5x2tcGH5N1
72E/L1+6A3OWhgFvmFcgFK8jzJkggGmyOT7TS3vGgfVOKYn46Zu6leCk1G5EyJuAvYENxWApVycj
A6Voi+/cpBMKEzQKRmLFE2titAvCcqkdaHME9xS+5HxQVLkVlF0fGWDgg601rByoqz8EdI398DuT
AXyJEFfEmhf3dEINBvekZzanbNAE6tWMW2eu63D+TGUPJdP4nIiT82KyUByizZXHA+2UiXPuXJX8
HiZM1osQg/+zRPGQ87G37MehPhCxZ82qM8pTzHmOEEjFStlL+ZycYb9VgZb6R01TZPlNUdavSVQb
rdbn20NmtDmIQ5uDBSCPKhiJW4bYLY4ftmLiKefCpSl+9mgCKdg32FesXErim5E+3W+4hLJep9Zj
6trKVPNRetXjJt4B6Ca8/6VZI1dasNfyNkDxiTTo5LymsWXp5gBAMMED00JedWuxQ27tEpmdL/39
yj+2wNBCOwEvCJiug5p7CEM7CsIYT/DkaLdcn+Y+9h/Ge86BABEY+yw0UvgI5FMcPmqAt+XPFuTx
+p5gpvEVNX/mjizbCObou7NRPT4XM4kK1fi9+RU5u9tW8o4ZCYQIF2WVUU7518mTcqc9JjLx2CBz
TJiEFLM1To6Xh4kgOcycTyKPeTwW68TfZHUQyxvxbg0eOaKOQHouNkbNx4n3GXWTON8BfRLuX97W
vOz64JWMLVoOfcOBy6brrTiTrOMjzFU/fEKWL3oDUUEF7p2rQHs5tT/dOIf05o4QR2LM496NtqjT
gL4WnIY1+vNuZkpM3AVfJb1A3DdlYFHfbPqags1c2iNjkqg6MGApTLDeDl9MQM4PN6MXz3i8kFX4
6PL17BLD4E2Wqx/+zf7E2wspZ31kwwbuVFiPyXQEJCZTDn2plKKKiF2NZN8hypEptP5a8FP71v/z
KAS/WvsP8WSbgO+5T0SzUS13I9bqlQWKTI70yVxvH8SpFVXtvTRci880bDInDqXpCK00/SndB+H3
ds59VDAWaQXRLpKqIKV93xLIjDAsy2OtDjK7lvSaggQ2jcQNfM70aYhvTw91De52VjW7musM4M99
tTktZaG7qisB/17Z1W1hy3DwuSniY1K5vClYIKACq3oydFY+6kk7OGJ1eu97wJMQOFbeTMRHnWvs
mBuNdZReIm03LfAFB2pvFwUlBlq8mJgbRLCXtwGARXO2vjoAKVkP9bqTpMxJ/JoCN7gew1eOObyw
um9shi2yh5YUd/zD7w0WyFlTYXcS0giNBcU534kTM6z5f91GWlizvKrNG8eCEX58P3CrkJMfv50M
0nqgPd/YAgH0CkJ0b+1VPA2GRSpASHBvycb9blSaCuVoYfFXMk/kDulbGWcMBi0QA2flUkLQBViH
ZVZ8yAu32EK93nL1VBp3sJ8Aleg+AZyLvsVmIQh+RbF3Vdn0d4IzZjt9cekZxm7uG7x3jxLoBKtp
ZjiEp/zRJOhO48a93YqIh7YjoIid8pSfDDzzLeCvbdGvEjzjjCJGYu/9LOkpXhiiqmLX7JCasoTf
jH+Qu5GXLd/Qw6LGg9iTk8saz0+K1dUmjmzgqcSUnLmvfVdVWh5Gfxw6peMy/AeuIqEPOA5XAsi4
7diLvelny1OJstcCF0/sTbxtqgD2T1qCjJ28uA/d4687fHhKiptTt1G9NxnzJ+0HhfUx42Pynopc
iUhhu/jIj6E1yXBNtgfhASdjf+UyoHCisxQTZMUWKtOLoCfdmzgS7OSbF9WDfuL0Six/fJu/q1bj
eru4LcBOK/oGzKd8KCaP2r7qjnWQAGnUA1U6j81mgoGSws6LXDQT/MxUALv6LXZhm+X+R+j7HwmB
FBBTWsp+ZgYAjJSy0lzVEE/G1TXT4NPqA5TPwYCZ7iLViZR/UmeY17MLBBBlRbOCRCEMAhAON/ca
SlZemgmLbyWl7FdTCmMyIbOXU4TwQqqUmgkZlIUfnbKAhkkWxu3GyaTpMwi3FmnX39ZbhUQeeasW
LSbZfhZPuqQRqYgt7++jdfeyOc4FU74Q/B+xVF0Cb71en21mmv+5HriTXcwWwOr1X8dMW3zB+nK5
taL3m7yAe6HHDOWrWdqYXNK0PmRNEhBlmlSJPVi5vgMvKPL2AL2dxZcf3vuwlkMcTPDRoezq2eNl
hLO7EnGdwNNGT6yflmocv8L/jTJtR6HZXd0YNzmqCSyLOqhGItwJf+NMV5oY/uB3+5bCeSPvZ3ee
F9heahaFZswIoYb8xTNYfQNU0M0VO1T4OdM5sv9kN1CtvDJe/+IuXTjKeOZDxuOS7rInT5ERqNRk
b9MihvA0Y3hOXAXrioq07F5D/r6AFjCCSp3yxp4dz7oqkMd4HyZl0mO1mH47eYmTisKlH3lLd4gj
TZhygYQ8e5PRAbIDpotDCdyJUIOGudNyNSiBjDA10sU6CEq29r5CPR6hqF8gv9Fop/IbhshhMy8N
a5QdZR5legYX7zKVYAK2wta/w//O3cJ1rVDLZ4ZHLIdZnUufAcKp4jKZDToX8lEb06+TP9SIpqxT
yUCFHqJ7nuLqRWxnkx40jh2Ev/di74g66Kgccjai8L3u73uFglGzxZ+qD5N+ZnwlNl/d2ot5/b23
UXWAz4/WDvD9jLWiweA+DVxJSlFpG6hbYvOhaevExmyQCfzN0v5ypluX4ld3vBP5oX4X9Gbu77TA
RUJR7mJzW+xoAwBC4KgI9NRTsls1nl0OKF0fKZYjsyyFJ1n5wA7QXN4orYRP8lZHJYRFS8UONuJs
pOknsFxTuKWZ9SHiC8TI1KRqJAtDS4yw9HJH41dxmpKpgyqlKg0TOUe5ZWX7V7UGuluR/WbGeT+8
ZPo9IHKr+HogJFmmYmaH1cXGgBWRVfOqX8Ezv0CxnPYejgrUY6cJZVKdZxnej69q3XLGrTyvi4nQ
3YsKIFPC4UhZuD+KFvOWJnIRC6ZgaANW22iMizHdFpFOD5PMYbMYStxFWwW6ByP4xdJQxbX9ZRDD
huVGXsAlSI+Omz/k/bLp5pnktVdBErS5KFZe01jC8q1HzU14BlZW7dIhjaesSb1R7oZhAFssAuY2
AfVULNpY5aOTdu3P1UKmoketF62b11SC5YTMC1ZlXTQ4TYvleIW26FRhxF8tHFWRqXU2ap5tXwGS
MIME4/Mz7Z5fyPW5kipijKvDLnpizqEg5tUy9npqfV72fEYnlNHsiNmnM6uHkSDKRA9rsceSsUr9
coRbACGw1srZ+/LpuZyjUQxGSJaawnZ/2QeZi34azCVwk2/yLY6ormqPCR3p2PjFKIMlgC4sv3XT
JqC0u6rV8Z9MZ7WSPd8GCA3BS/ojF21czMpMTqIe+9Kd5kbwOiMDZPpUfSwycG9JN7Kbjn8XuHfD
BN3nUsycY+whAPR+5wilZF4Qb/oRmyUd6CmJ8zbSkAi6aczLZsC6dkB9UFpC/l4kBInADMnIsRBa
Ogtpibw0XipSVgkYILCQOoVzdWsP8fhA2Gvk7EY0BpFFJoedAXqdMNZ6dUXl2Dj/w8YtkWKnlNqo
41nwMz5bYF+Pa09ZrADE30Jlc9VutrBGgWd/MbwtOG6pzxH/gEg9QhC4lLlOsDU1hjPm+paavAYD
3OkeQ/TeaXnYTkmVq2Njix+NR71rvzCWAZsGjtCm0x3uJOLyM7Mj8cm6ibbe9uzgSuiCleAvMCoo
2tZI6xtfTiN3QHIY7VJrEAqz0EI/VTwB+HxtYDVxQGbCIy/RCgB6ORQUSvZQrGam7tML5nIj9iLQ
LqCOwUohTTZ9b/rp7QpAHSTN01hgALHUBTrjIAUrKzQuQVKTSR8SL/NAbUeMf/GAhas7RjG5ZDJg
ycl2I8a9VkkFLE5ocNJdFoW+vCgirqTLJLDSemgrTyMMpJM96oZMFS/eoCQAVOrXxnFppRkQntdf
bELC+bWaZysdzAKWfdKrkffyeEHwJr8HLlqVCOuTuKGtyMb9TW3NwePsHKGLn3IwnRyO9Y84yxzD
1Qzg7RxLo+87oKCh5dcFMlTDtuWgV1NqzuylzQY7kfgIoeWLrT2uWnd9rRRYI2F2wvK+6+AESp2p
qSsWeYrev1UYvJKVjNBYohYNEIMQoWCgbNAD6uAp8A0/JDV3mCLVZQLsPMWZPAhwNu0dwcdzBviW
5vIm3zGiHemXfBlOKFo+oteHdu4axNbev1/RYVrzLa5y9W6Pc5Z+R/jt3G58bjCIWtvKljhZUHXO
hR6rn2sEmBzdvi1XbtfAQ0OvzW5VMK91F5pUIVtYT9VVkhFSgwdnWxzDTiG/ismKy/wtMCJtmB9v
DfXbyNGHJcnNf11HkC+EXcBEuOen0aqh33Wcef7OnG29wMIW3iftMps//mvVsbZgXvq30rOUob3M
PoR0U7QRcN1VHke0Pu6aThYtBn5WUJaBCrxWUNJFg7gh49B+nBmae76XKsJV8OYLshreG2uQdVFh
1a3/LbrpIYar3gc82Vi1R+CnYkCq3W8cevSEfOFlVxp64o6xMB2pDF1VeoX82YmrzuNtQCZNDWTS
tW7NGjdwUltref5bqP3wV8yzAXltoea3+kki+RHVg3oQ8Ua5pL+s3pwMrKtTMsGJEaWahWqmdlCd
sKCDqJ+gEeokZ0ZDAuhHsPaAJlFZowopOwo4Jbzrkm4OCQI7wv5n81YRC/7KkxzYY24SJ5diSAce
jDOKMn2kTUMo3HaYxcF+oenAK20Ug2ia8VY/gOXqglxCkJgu5B65463xuUttH3MQ8FoGCfqlwaDH
QfaLAi7+pD6Snx/GPN0HV2t8rFetBDnuRcT3D8VV/fQKcq+TpByipnido2LN6cl/PSmXYXpY+rJs
wJwjODhLxrTRWLuAXCa+PAzAcNu609UPJe69RXOmLvwNhz6GpEUk0i5c7qdhNxiJZS0rT47pi37l
yE/Mzq2JpcvP8VhbB1HuZPp0wEFqnwoZudwVAeriL74FaFSwikvJVA+9thUK3ldvGJuMj7XsllFF
p799atVJtGl7ZnDd7Tv3CYye0NMG6NTOJ5AWwtRR6ovLVLdo+LsMYfOUQ99qhT+4xQimBY95iaDT
bnCFA/5LO/01bUR31f4ECR2TReKs1MK1kEE9aZICvnwt3oBbfP4ylDyDYcr+WsTLEEPJHZ+0VNCq
POSScbMIdLS9qu4MeGNBilEi8+5/FIc/vh/on6ytcDUae20ozz3BR+GVdxBjkAB+C8DD9POsfiIT
lF3bl5h9Ql3m9D+lNum1jQTbHS41tILqgmDKuKdf9fgzqfGuf/lPbQJ39VN+wbZQK75oXnJM17HL
l1YNbuJyNc89un4BPYvCFeyq8f+r7JtLjzSiZguw4Wk7Mf7RWKd0JVlw3fHzMihvaojTxPtiNpq7
S2gV24NtklAFZDZYJFdrE+s8D3rCZq8JmBAO0DD38m4vC3Bbzrp5nG8E+dOLptBt3qP/gGBdneOD
t3tB4pf1MWlNdLoQLvmKVLsdlTCilclmIEugj6sOJl4Fzhwm5yylEf1BuP4nNY7JlM5LlBmzqnBI
HNIPdARAaCaDU1aRM5HPMgZ4okzCprWSHxzAy0dt7RbltFEb/HzDwnPXGBX+fU4rdrosQHvBjreX
qPFGVcwxvkudk9gfIna4l4cc3WGckAO5Ek9UXCNGREfir00ZB3iOC8t1B14W2DNTaA0Fi9Gp8fTY
qJd8vmDxuhk+fb6lKrjRB7WdPFthtoe3L3hUaZKAZVE2W15pIbo2x40iZZTIXq5DtSetOXs0QIWb
497ea6dp4N4XC9jogH92k8dKcL4eV9+sxQItG7OfztFPJBVoSGDNWH0+xJkCafT6gCq8P6jT1Fp8
mDUNbnBg+Fp+vI2CuHbDoZXdZuv2rZaTFwprS6MSftHgJj5aswdw3EDaebM2iAT+IIP3cPkhB2vD
aYZd0J5y5VCKeyxNjpnYuXszcIlJiKXhC7ZNRwf/njQi6B+Ioq47HalljDqOr//xP75g2hFZAcGY
lAzbGUVLmYg2Leeyh1BJNMPfbDORRLMBKZA+ptKh4jAaH2CozsP9cIZkjyYVUZWwX2AcFOOQCW1U
AxcetVTzb9X8KSmZGB9SBLu6seOJr18zFu8GSn+kMIxfsH7bxbi+sd+clGnXNyvMhmflNXSQTZpz
t/WB24/rutzZs8OqGfGkmQfhJWJhAaPTFrjBe68CDgsiwyBK/1kxfZyKzOsR0KgIj5Hxn+HWVc59
u2XSBnTh3vC29gojqKMKZ6BOsIQDSBOfllG0CbFWUwQRqwhMOtKYQTQguS5MHVVpOA7tI9Z5M7pI
kSbydXGHh7bnRh3Ns501HWwyWI35xo+qmj/nijgmBjpQojxkg27zNDSY4BEYKe9LClz8ipqKR0zE
0J0GTzh+EYrAB8asphoCdrhxFeuJQJ4QaZU2YTXSKv8XT8tsjpNcf4vJVuDLfTQVQP2Z1UzIt+I8
Dl45NluAmh2PlgnIlw50PF2sZuxAzIAOtsquEixPGcvHQBdLw3vOyyPlbd3zDdPM1Dgtabnaw8nt
REbk9lAW5iFGjIqQ6wv5T24ekxfYQRufMH8I01gTbhs1DPbpPo0/JBnISy9rO7N2noEyNCCz2KLY
lQLt5nCMCHd5mq6+rqYtIateR7gC31hkZXqZmWreU2fABJ3Sdg3b2JjR5oCznonMAaooKGNlGBWW
YHrVQRjW3eutO9PrAkW6xFiRYmuXLVHaWsLl0XheCBpfoWM4CRuH0QqYTOiOJPf6og3v7v5HMQjH
ySa5hB8VvfIxtruc8nxMhERhbleAx50xJB5GgZ7mZ5cjddPoP9F9Z5LenxGh9GhXKHkmQFjvpP/i
L5m4w50Bj9HOjXdkCBiqN6RAPbEbUOo0oRSj/1WTpTVDqSNxabLRiOook8fJ/jiKeYciBWPCX/Ho
xjCH110BGkjvO4JU1Z2+drV63tbtB7/QSJN4HHE9mgT51hTZIhmutjDrTW8zC93ALXtZGCZkfOLy
yJG6vlqep31eUlWiXeovuIV53fMTRKOdE0w+N2Tj7jJzbvBZix5H/L9tFEsfttWBNW3NIKMVyVuc
h2aqakKI2FUsb3GCe4/RBE2L4hKFnz4X4cY4OYW8HB6KfqeKJtvBgNJ9w/tf8WQrdrUHj8VyP+Rj
EMY+w0cMP05lGX+pRXKwRLlG00q9vzfqnzv+jKFN3E9HeYxKLQp8g6xy9FXxxGAIHynaRvvrffgk
UvK1yQBdIYoSHIJkJd5iMTDKw1Qv3eMdG0cBizEWYEocrZ3ZFcOQTf0nK1n7FsoQu4idEEr1Q4VI
rE9bsQ7aDVHzRVBkWiMb/Tm1IYMFWkC3F8dV2+MpzZ3ex/0+zbfr5gz02ozXD47Vaqi1IU7hKzch
5ffr4Z4OFCxYqFvet16sPMzQSTJGUpUm2+gpURJcXBFGhwW+3PXrZY3EXKBez60vsyQZdbj1uurU
Q8kxXNbTAUmWpma945qBpfJbE1xY61xjy4ocO99fEIsxiU+NsJqM75XiYGNrQVGrLhn8HP+OlMPX
D/EXXLVn/jIT977F+pp7ApBbjLhRo/mhdIn9NWyZMwn5RS6UGpoq7sY7oCrr3AdlT0970RHhiYt7
eVhv2PL+1RzHMhIAieSWizPZrFEjgmisFf/WVAqKd9N7WFZZ8HPThs8g4nFcbmzWTjBm8P8E0syn
fxxELcTVf2aL5gZw0sZW//aKrlbCMQuQgWR3xhNKmyeMQATmYD97nKDPCPk7so2c6OxQPNiOdiIb
YmkpP96Xyux45aLWvHRTpEz9xbUlEYdKKvuk2n/870Qx81MX4OvIq/V1+B1J7e+yaXbDJJed36wJ
8qmsWJFoQgFk6xlatKvSouIJOGwTKJ4zaeYmu6msewrT0tD6h70nziTUeBRHhkKQ4wdGXf4Ub7An
YH+j/KmFY+3Oi1COQYem1xejDvyBuYb1Bpp+lPPcJmr1k79RwA4DYruALsAmhcFPae6OAb7BShC1
OY8FcItvbkshvDY1lRCXuxPxDe6UF4aDO0ulB3a4ke1oCAXE6wCi87IGSjpB8/e1c4ZQgdGda4Co
6N1zqkivabpmJzr1+IoPELI950vviYydgMLkRK1JfRJuauuijdOxQOnRsxWS+P3UZBxtqG798Y0y
NdqgxagYt7EsSvLHuql+WEFEbpovc2pc5eq7O9eJLG3CGC/MW4zeaN0Wfg60HvA9jTpwlhll5hX0
KynOZ6njuNXejdgXXfH74fXwlis9347qqp0FOHl1xTmwgUaTs8HDJsHMknoc0osfgvXDfk3y1zC5
eRGl8Em2OIF6/XMvdPF9tbGWbDdjEFiZXQKjQEwnecxlJsLkEZGf+NYf1F9i/w/nk9EIPnqkoFRB
Ca/uNRvrT6rOCASEvw+83WEiCtaiZqV7JbWe291fcOiXapqhPkCih3eU0pYcfVyjkoexZWU/8F4v
PMcz5oks3Ny5vxRBsZeeTkfR4OE5Jcw5IG6g0G3l3iIDa2Bt2/pdlmi6lKyCVnS2VvO7FQXl2x4/
1vSK/ty5jn/0IVybQwOQLCyj1s+UNy62q69aXQfPxgH6rxjsEvHxtCyEU12R6XEeajHBZsDbpTqv
cCspnnXbok/f3da68eIxoko3/XpTo619a9d6XPLG1QrDO2yw3/d/LZ9+0suD7GY5sdz5ddtiM179
clvTMtrjSHCDfkpwkdU4PK1CPoKJA6nEOvMACw2RN1urcpA53Erwn8UAks/4VUzFSRbiOyGA2fbU
ACL09MlS83oSz7/OYXTBgKMP909e3dDXrj8+My63N1xmoYZ2m23gD4VIgBtv1xlzg2GMV5PCqE67
OIPA6rEeLck7IA0Lipa3JW6jD0zoESXRoOI4XsZSimE5j43ENtYjdVKCK7wsVYhYbbdxQptSGsHl
12QaggNhLEIy4d8Z3E+V8IhIhqlCar1RBLJ9Y+23kEMbydirjnP05EW3TIAoiBTq0XZ3cVGe6j2m
BgE8VpKTaHxNr7wisSxY+8CiY1M5pDX32hqcIFqz33gAV/rKAWdL89O7L3qGOqC3mW7vG9bnFtkp
j3nXUIC8cpZ3aB+n+Iq+ImmytA2OiR3lcsbYpRXz3ZdINom5znblNshHQRjXT1Y3tzlCKtYcGmG5
9p2APduaxEeNJZzCwBSdVLguRvT2ibQd++EBmEcydyaAIsiQ/q6GA+lDZLPEOwsHGEDhKioaPGDY
r+CoaTc2IIWwA8u6cbKbp7Oh8AYGyQ5JzYpkS/aWFGhDsNDhbkbxnXV4ee3T5MC0OKSqNEEuCSVR
CF9AHEw8mJwvzmJfOpOr7QjJtuoUjWxi+fx+PJBXVhhyOXd7Rkv/ak9XQ6cTapId4Yeoo593IN6U
aEIM/EtAB3j7bN5b6W8+wp3tirV9FIOhTe76K/3vTZNauALADP10dIJwIhBUf74MzHgvXaubCma4
ZzMU80MHR6mzwnYgEIV9p4omcU7jrpTwpaS9+EWUhsY5ZXVSx6sXRMUZ8vil8R+sMTF8T2hF53Ig
gXgPdgKsP3dRD7OgigYh1PLmQe7w+ysSJ9hYVc3ud/j4YihXboOUcO13I+SOXIOXCqif/bNFxAZM
R6CsTUpLv/5xUHe0R1KFR1OK4KE03Jwi9f0HdiOMVfRK5imPa5qKj1NOJ3kwGXXZ1n3f7J7p8oSw
ny0pOHioKXBO9oejZYaegTYzZdLbeXIjM3HSDcY8qzN+J9nkLaBJKWx3e5pxWsCs+9efr1sjmE0G
/Sa6OvJT1ZzkLPeaKKbK748yiSauLzoLtiXXUM9EA15PoPnqE2X9CdzvvHL99zomydcLuLDPlJyV
b0DnYZLCEvNMgR7bWLDkWkdFc1ZYRmrMbYDrz/xctErbzH69fi/970VIglUQpK1zM0rHhBUi5wn1
p1DhB4Ab5fwsC24Q2XN944FFKusQexqczhtFjWXN66WA/l6MlkAF0Gn80wdwCBSg8lafmcR1GQtC
mFRoC3Jnno9m4o8kvsfeC8HR/LSqARiFbMmhQts+f3HwtxzgfDQSyOS5Zyi/nqg/UMMrv6ZO/R4c
B+tiZkjxD47B6cJyrP3SksIM1lQbZFJWS3xYsWxZMz777fGLYKXr0sYB2WMyAruk6LNHxbxDUT0D
Ry9Ahsfru2gXAFpUm74nYpEA3q3xJTlqtxY8+peJ7WhWTW/VNcBrKNPw/DCGepYh70WnlwISeR+E
oD8sJAfbJPPNz7VBmCh/dUoeWJqfxgKyf+JwxQ8k8/cbb4+YpWQPV6rLi4MlSEf7Hko+LMjC67GS
T8NcYzPXdK242/X0tJBXnCSdpHJ3fARsbi4rYp2haCjoG5IuKam+1qsqacveaY953Kbs7ZvCeZhe
MLudiscGsxO8ZqTEfydSFkyPk8IbSApGI0fzc4q3vnVv2GPoRpbyeChAliDTLC1uhuqOtl1aiL7s
R3aP3aafpSinbWVQ08YfbqNev/w9CL3uuYrpoUB1un6yIW+thfo1UdQnqtdDo+x1j9x/jpX6sV/Q
J1qieN6Tu74uyBpfQWFydZYiVVwDb5tojZb3wnW81r17EJTiQb9Tel0KNy+TiYxlxM/Tmx9RkN13
ENgl2c/kAx7AgfPMi2Ij5coRsv7E8noat8jZsuUckvAhuNdCE5l8u5HdHmm/dAMxo/HywSUxCrJ4
TQM8TQePDx3Fez1tBo/YNoQnFnfYQnyDdOkjvHC0BHTQuWZP0rHTOgjB2VG+wRGMTKhtf0+EqB0k
ktDqhYPLYjfuobHMnWS+LigmUUBzIkYmIQ4zLur91ftTcemhw0BnWjdcLxodngvTaiNM0u1luH0s
NI1b1qgsNsOJixcJyEDgpKjWtvbZJrmiVjm5YMmcEb1ANQhqljE7ywJzTV39fO9KWO+bUvv1Eo7Y
PIZW56szqdnzf63UaQIwdu74G0yHuQ4LYyM53sMwSjjWTezni1njdly7/PN1PmDhLICFwIww82Rg
78kPMh7VElnSJ7HJlRPNZf9jBUpicCRPgYPF6qs7BNV+nOz2zKsTib3cyhl51vRRqvDU06/qauGz
fV9KO3Ji0qylfuHGFbv/Hq76gbhKCZocOTswNq6N63wrgABxpWnii9afLQcUddbSpVD+ALqoXyF3
s0TJifKol2Hof9qQuPtkieNXNLvPN8Os7sXY8UJi9bwunZYdOjaTDIAGesHgJYM7o9HiYua2gG2U
clH1e5Otl/WrQwEczch77ITfiOvQw+e5T3yeTxvgs0KIdVRjzgS0aIN1a6ONwVf1KM9JmeAUJWUI
LBmD4tHdxNKnFOVvNGHZzjfdgRxm8RurJZFLCZ6jDd5+oIMKHEZdE5hhGPHOYlZfmBsSB46QbZk7
VN0Gkcrg7N//zUs2/KJ1F97BEzL1gpY7BoW8ZY425pJvNm2HGbEO6iP54VOFVIX54eowWBg6z4J3
JOxgRfZMqfa+RjEgAQpbkFrN5xAndFJDpP2um9nzv2IOxDQDmkKZYahzcA9L2meWOsKP2n2bmvBQ
467QoUP2LadX9RQ76KqOHw1aSmixC+8Qo/xcllAAGVIMTpLG8a2bzfSaiAxZ1/zhWwUEbPGtKo6C
ls93UN2lnHOWmeen8i7vmM9S49wabSAFuUlWFKRttjMiDdgqGDHQh9NuA8g6sqt3K7P5x0UopW8p
GvGDKKrdxoqgXC0RVQ6n79pPONj2BSenk5cZNmYPEg13X1JtllyuT+KNsS81Z7EOYug+GYBiuV04
XoXiBIryumSf+GUX4qIhzbG8aYXcLqd62vCFc08a3tkNgQ5CdXTZxH19hCc1qaqxP+8UIoFOLFjL
VYY3dYeMJS6ojuSoXcHrjhPrU0uYEwBup7D5pyOpp02iC4eUJs8k4iZ5TV/4Nchq0E15ZLBXznPZ
09M31NFGmFHIF1WhXTIN7e4suqvUjAcF0mG5iWaoG3xx7LwWi8gpB8CDo5QdTZnMYJhkBV0OCHqg
pf+i7eYoDnuyqw1gmi8WifNk30JHRfIL4baLSOgQWAF7zVxzCheol5aRVZuBECnqdYCgn5Ne8VS1
jHFGbsmB9+TKLhWYiLDdeBJjsY7o0R9gq9iv4JtnPd/Aic2sc9I3OMXtZ7mqmD5tnbo1qr+wCsJP
eKO1IhTzHXIRhU7B5WBCLlj766NYMHsmrqmjF+mL9H/BDM8Xky4fwIFtHQ3hqX0NBspoOD0Q0D5Y
4u7EvjUOxq9NPdQDM3tHxAKYriutBEjt9VY2qMbrLyX8zCbXwp5fQoB0pFB2NRuKaDVSHLsy4FQz
vXi9vlvYBZc3F8bEiOUtmX+0vKqCiNJQ+Zd2WFEMUsQKFJuLU/+qfQjF/j/k+VMTq6UrbaVb12wK
aBxNq9LQqfjLpgbqFq4K6hVNmXOyFrJGhhU41VSS9veNnOq+L42pNCsxiQoa4xeAdlZSuDQN+6jT
ti+6gzYsmO8MEBhJMamo7yWGf7SJ9tHBr6TifQ7eart55RaLy66IxHYP/UVvvVAO1VF9gozyzQ3Y
wBS1cBIwKZZLayVLY9FSV5/+LBLmMyf+N1vA5mx28oW3R9ZHE3Od+F0XhIuWlOlJw3ICMyabjVUm
RpJEy5pHhlAjckGrQrkf8oFwa5Lh1QLA+ckg2lH/Ifoao6Cv26sRu800ruoy1UQCHP5kezW+ngQo
yIpqszoo5m7ca1PmU+vwxk5ttRRZ4pthmnXbijHFp9gIZ+/1jKhe20GIRpHK3+uYiehVWX3ZUJ3R
dUhHBFryTJYuV2P7nMSLjG7OwQwRUirrmg0oZRitA1XlBKCZSPO9zpNgO+qISZIVqJbSaT+M7IIG
5J0Zb4bwKyojFJno79ThcV8tnGKEvR6ZZ7PXsBs92vYzJBwO8spdx4iSDnF4LIhLFAVTofm93JUW
2rBTXGZt0VXMu47t38ulzlYK6vnnXopB46oCj8RKpHH7HnLG5zLyk28xriT/gfKMbW4C1ADPTSDn
QdiDZarwbs+1DU2xLwttXqwyQljPRfI2OOsf1Ix2bZUQq+bkuTC0NWo1sZ0AAE8IS5PZCc7sMLNc
Vfg+wz9M02+5XloxSlHoYjmWR9Nn9q4GgoVcIuPxmzxWFbAlUUSBRFxM0PcZMg/KmST0ll5lg9D1
xd/cE3GALOhGoLuixtFs+OqhPzQ6DRsFPn0SK/vmTR5VAr/YESbXrjC62vulyhay/szZMIfNt+ri
OA6nvVpG54x2M8YF7NeTxqS3GXOtwKRAoTM9d0D1cOWiDl4uSFHmF8kPt897LAbwmjvw616lc1ct
NwD+AMrEAJ7Nw+2ZLHr2mx+kfjIlgDPwUn4A4LmYSxlhx7vggPt7Yn9UyI038v4VBnkT5f444HfZ
fUOhd6V9PzhACWeKSnehi2ae/lQXZfkaLsYGInnX5GfTxNgu08JIIVNwY5ZyrmbjMSe7B3hqtYt7
tCj4U8yuK67Kvuo5W1TAJXMhLitWCYl1sxdG4yNbXZ1WyoE/DXfJlw3b7AkR4t2AAwR4v2RDON+H
PPK4/y0LbtHlEHV6Zr8j1lR180TwEh9bVFqE6YzllP4CePbJpenJkPkeMxklJAMv3/bPQdYZlt4s
92WSi51MSd91hD5iUYCacI96FczgXdXFSwBnvIjMrpJBeIGfvREAMTlsg/0Tg9tKeW5A6pxwnr60
uv2UCXzj5/dH2rL8MOvv/063akUFUo2M5GXtOxF2ClwO2E5mq34fqoB3u2aadMB5PsCS29sNH6Wr
sOReY1cYfvHp71gfPAi+m0hXPYXP63YxyLn/SIkKB95C86PcXqy1urbEePwEHkCkDOBPngkzyvGn
0R5uyoAqBXHDIbJflM0WYRrcToGhAdG0tIiu4r0SreYYqU0LY1mnzTensyCxEJ7dF4kCO6X3Vh/X
K7C915asm4Fg4SzQclF5IMawund/U+fjL9kTnaD2M7tgIkSn4ZZItxJJ5y3cryx+sq8/Wd4tIy5T
fLbcYrBOmJOO6Ds+wKlgSdZ8i4XzFHeFjkOOeHE8VrAJnc81JID6y23eS0uIwzzEe+vTifwKuxvY
IFDw4NjrhO4SLSVBLh+sXXgmmY/egqVCOz3bNUNd5+GOLJySDzFViZlHaSdSjlbyUej9y3yh8Dh/
Fv+aOWvQ3rvCROpaXcYujp1HOdW1N3xdUuIo3I8zYZqrp6SpvfJuWJHXMuomiAU+G+wJ8GCOt813
BfjXbxVvvBxDhojMYvaz1CcOb8d7jQDhrJa676F9Nyy6Po0GToqtTACJV+7m8TdXNc03eXKCI0qj
1vKIk0k/f3ERVctAlS5T+2UyPW0TzV2WSa3UYMpto2iD6lS1uVg5VcxU9uJgDW3WkYZfXpbq1N20
RA/isIqjHa1bd61E3zAJGWE/vz0sL8+N4JFqTOPxZGVNHMmwVisS1p1Enbgd/D1fYIY6tG+YVVrA
pBN9YYb5Lfl28mX5RdlNAi0LcKQDuhxWh5dmXYZlDOl9rr4FiHU0fmcCS8wS6uaUWaE/1p6Qd10l
73P81Nm8QW7zP8YD2EDDOvM2pMWlOK8+lWdDNmj+4CDALDbUka2yDJmM0e8emozuN8VxvWOvOBRs
Gyjvs9IxxNcwSyetwJ4Ojnpoeswgc14cBc8750nwcm9J/rFbD0TAvq2v1dP4Mf1rqB5utMDA2VU2
OG/m3+OqIOxhF/qB0koPipOuUHQsUAJ9BmJsEblQC06aJEMlq1WkFWDYVYeXiJg7Gj8S9zbqpmIW
Ek7rVMi801uMD03St1khWMT/vAXTORnnFW53SkeY8uUSA7HB+GLACLBqsEFyesoho+lkr09iVsy8
wrRjTjStfKIztCxd3F7lE+1oIY4f0IR7AVcIeK7wV+3bWOudNQRHbozQ0YxZyu4ANNDUyi0uQD26
pxLo7bZwyE2LdlVqY6e/EcaZpJvHJX+JCJ3Hxb7U/aghL0LAVRLxSLKUYl69yF5XcDkdYQSptXd6
rmPjf/NYibb2t9DRRkZc7/UwBw2EmaGtcYQa6wL66YDynp4sJ83H7QRbWLBd2syEiRGB3fYJ09ST
sICokBURwLegILzic2O290Hlvo5YbivyCTjaI0RmwVInCZYwtdUl4FvOdPgol37DF7VV6i0eLVhh
3+m2J4O3YGJaVmJKC1MUfByHIMLbu6nST8f6R+//bfAttjWtBtLd5K+1L3FEBwZ1588L19+YlOH6
UEwgoqzrWWNdNpNlhwBFPQpS4tqrCVfImBvrIWg87x0aNhYy5ulevCzEZw5Gy+eiC2JWNLHnchsx
Nu8S/sWKgypvd0p72bjw0/iPX3wXt84r5SVFVauwxucVwzyAZ791u5pBqNSwi8MeV1BN/5czbNju
+j079vFK6BBvsfhKsvX2kGKA0RYUYqjLi1Qpwm9KngoG78B8dPhKDE4xi4yFfd4n+3qUPnzHUQ0G
7ftR/5xxJGhhIkBAnKKs5TKznagXqUqYUeHpPpswXW9DQTjG3ARnjdmhNNzqgjdqpyL+aX0mxxG8
+PCBRSXPWBFnlLuSe/yKMNCI6YN4vIXmjTNLh65fSQgLnO4a9GUPG2f47+Hae8Hr7J8YO5NvN0e2
yal72uydYL303XqGkMbKw89K+kGYAgtDKdv0JYt1aUPzft1W0Vt2UnuNf/eEjzUCULh6WwBmDAt1
n+rty962V8V8U+uDyoGebDySx1hYttmsFgwaFAlb4OGuSGD6BcvDbvFEuajH4tyV37neaNoDgs2U
TSyuD0hi6NmKEEfFJmGwIIIQIq/2T0FEMfU6dmvchLWZH1JO6KHtf6AtO4nlgCp3wyEFJYd87ivR
IMD6tVewcoVul7rc/xKiZjPAJb6PKBGvX/EVIzU8r5gRx7DJDnlQuZVRhHvGkeFUN5IigIdS6j6s
fMJuxveUpAzOJTKC2nuIHMZGRfOBJQUMke5BnrK5LoI+OeivSvmLKQPEh4EMtVp/3wMqu+BMa0Wa
GuMM94fd7zxmBm9oVcbPFN+5ymB/CBuoVKmWDqKPTbt5lgP8C0fdL7IM6KSh1P5wjkQ6VtlKQIxb
YXUg+AaH9k+o8ltJ+1Mf9buoY5UYpzhLhQrnLu5Tg5eTSkxIrRC+hAqDNZsernAuC0M3p31QYaRi
Ohr+QDodWKzn9d8zK3VDucOyMKdbzVxg82WsC2hoRsx19cwJoh8uLjJOqMBYQm8G87JgujlXRk0w
aTCwrF0cS4Gc/f9jMNx0aiKN87f1L45V92BengyN+NPBuO4x/1VV2DiRXov3MMBA9igQSnjSAHy7
R3/uSeZFjgY4oRrkWBVGTMZ5FprdcnxLTGlGBM0+QnKinBiRVPoIMgI/12o2b0PI3QUsVzU7sHb9
P4A2yD4KW/3EIJv5Ykrfrmuv4EzyiNaRc59vcrkm+8vDo9ERuK3JyHElYCvFrraXOkdf5aq+yXoC
N5GoA88FykuKW/H/SwyKTTSo0m1ecSscaafKkII1ii2LWFjhjCT2VsPgnTY+aSb7pPcGYva+7gX6
JjmbWkAZW3TK3KIZbG8XlIwPi609mQLrUr6kSog14UUPLZYss9+zgyZebUaglNxv/vLQhfYX0CQE
SIEhTVKkS5a+kRm6W0lZKBLzr7SWHiPh9v/ynkeUXaQgAwEzebHI/gXCs7oG2lSwnIb4e9AqXCJ6
DLm9nKQDho4VfAMfeNYl15BpPDcxLAHF8CCltULf8NkWJRWIq8P0nEqKyRz5UinpJdLdqZbf+s2i
JZejnJEmXAxaf2bnDnmQI9LLGJkOi1LB1egnfgm/Iuj/7o3pEnByQErT+ImgCi8j0sBGc6hSP7hG
WBUoZPtT+kI/h22Y4PYvv8CDCpYrKovQXuiu78A60ceJlHbogiAGjeywluqOBMXQeVNYvErvf6pd
6Zb5833vkYEXDuFXQ/vDzjYcUJiPLnUi2VWyIZVM/zvCfETb3+lsu3xaR73jr7BvwoQwYNV9XFta
vp9AyDrd/QO1oRYGCOxof6LGop5xUOQg3cHA328ZBO1xyYOrFhTFVXHdd21amLl3twWit5Ar2/2e
NTKOA3D6hk+7A+d61PBKjUzGZCNwEYKF9z8DcZXTicxSrSEryi2hM8nKCdyXs2aLO4gPHPlZ5GQf
ko4nfBRhf5absdNu1EO4jQoEjsGAZmUYUjQw5bI+qxNM4qlW6lHPjdfTRd6uFTGwmLUF+lVsfix5
vmGELwsUa8/rsQCIpL7zpxBrVfOzbJZKMp/O665vxbGrIkCvnW0BzkEtEvtLtcKWg0m7uZsC5KsP
pDMcugjHhuWw1HYaNG2sENU8EkIDsck4683NfM7EV08eNWJWeem8KEcaRYXNrB74ecne4bUoE3kc
srq3yqezyKnrOZgEfspyn7SzY8QIwjpPqFbtf03o+U/7kfmDJtZkONySRPRw+Z1F/1R0+UtGyufx
zBeIQSvanUxTK4auZSkXHjG2bHqMgBa3zTPpfdy4NjGmxbc7bEqvrE4PvGFbBa3bePv8UfyUyOdv
4TJWm4IZZc2a9DUHcLoplGzPQgIUYgeqJScf+Z57M83Ow3I6Sot8VHHN73n+/x/LMhCtsmgXIPeJ
H+MzNDHHYMSNmhx6zPm9LFLmDBeqgRe58n3ExjNwU1tUlhOGqD1PVniTmqTeA6Zu1G6iGBpF/4lm
3a9lp7rYGv4mAWnhChTESU9hiJ3RtU5e8RXsP6oQXLXj59DNk50yCaockGPB+cpScghOGNCE9zik
kz2w3Yo2SiXqdqeP2XrfL67vnPNs0V4pCCMcUtdLSAYpGM/UmNZ5SsKaEorygB9KJ1YO8Sq8llID
fu66QHcvF/BsvqDBEceli61bMoHfShcr+OAUINwxw636ipzQnsUOyDvymOTyb2lNXZ1kIMyXnAY7
kjglYbw/oNmQDZUIuwIYlzN8XpmXRqGrfvdLMvbJCGZEO7ZKaCl938SVQY3GqB5yyRf+2iZqWBmp
p+lrOl/8+HAoeE42c6u5JqhQ7galdjXt7cQHxP/ss60PKnVJUgAt1W65fGD42hFCD9N6b1Sc6Yqd
gXpiLvVmue6g/IhfhR6mbZ21YBPWyC4NCSJstt5LNF8Jz98bk+Gw/UDIMG5alb3P2VBNsave0/WH
4gWLR9riqScpCArGzgs1MouW/6yyGG4WNkBsVjOspM6ROAwTm7Y6+9vd2TnBi/6GHM2grNQnvXO1
h7/1MigaKtJlXhBNirzuGsykLgz1TDMktiTNus/qcnBDaXLD+3MGlUYcmRm1/Acvj0p8DdvAF5sI
f0cirX6jJOaN9afiIkwOq0/tHnsmaR3o5aG1rkUWDxUkq4tb97j9jmyFzJxbbEYSRYRGEHmjVzyk
4XV105nFFCZXrhD9ZsthaCZk8MqqNujW720aIIcyO3kY7NXEDNyysdHsZ/bZL2Obq/ZXtq/Pkkyr
+s+JSzIbashsY5Eo8hqXTwmjZ24OUWKGCVRslylwDmFOqLhw77Hqsi7nqW074gurdjdmCqEWz1hB
3g5rK6U+hRusc/h0wspjFOuCIYVH0Amq5xFoTlPmbG0RV+EsIiDXpU0WF+Vc7qp4g06fDBPqnueK
JziuOUOBYzmFTTlNG2r3ymAPbpQBM+d662cZDQBLlWikgdjXIx0TIUbE5EtnXAjY9UN7zxB7QlJ0
31ovanJ5z+SE3F/9JW5KlmY0wuIKnJeIFn1oLrbVo0dL6ts7MV32OBYe0UxpjN+WyOlXoNGh/79c
x9kh9oYAjUNVBi5SGDk2dheju7wyapfzcmjnQGZXVUeU1/X8ii62XWtYKQpsznz1bcsLfj97UZNF
qIl6vYudiVj7kHO5Fze+ZclRAG60TO8rPdg1yfG7B7gmTNHoD7Kkpw98emmug4sWo0j54OhPOtLK
PCZL8pQlyxrk8evjcF/AqdUDpd9Ix7JdQENyUL8M+kNZr7iQJn+jHATGxFR9ZxgwahgRxsonUg1g
P7dhcfT8FzgqvvYuYGiEI1O4fiOrhHdRPioTCrEAfTXbVylMpzdKGXfhgU/siiiRY8mMJ9nrskVN
DZqLx825gEsAD0Ado54egfFMXob1+SlrWwu1GdGdgs10FO5h5jsCYlQdOowmyhJHv4eI5go6q3lp
Pz7T2ca+shC1x4aWbtqEyJCKf1OLueQNIqtEPPoh9gmVbk3Q17nAUB39lwomDPgwDXtXdStW2OT1
ODtJp63a19KOMVcAXZ6wQ5NWPT6JMybk1PppHV6RhbZH5fb6sVrVke6Zp3Tws2p2lIOmW7QSIGmi
clS+IUtJHifoLEiJ8Es9mx3M/SQmLK4SDin0PoTaomkdQlamCUezdkZpKcq1+uPAllqf79KlU4el
AE9jBN3XryPNeKEP7etEAqelDXuwaJgsjpeK+1bDW3bvI/w11bzY8JrcaaYK51jqzl/uXD+82PG8
fPv89cFWoV6VlX5hCF2e4/H/dbz/9qNkE+hWZXxJfxLklFjhmBqFE83t4T5EA0rVJ7j7304GYQz7
Y503xwF0xdimdgj3boHhP5y4knB6ZvTZE/KIemC9zlHmF22tpIaMy9jCWinODN1HRjiGRtYf1i7o
AJPqEXlRYa0VWXi1Zood8C5JQZ+qvaogMwBuiC8maICBQNylm8/ft6PUkZBYRDNRAAiZURMLhYUd
Q1HLs6CT9pzBM7C9iAhOofeqSI4LrPXjCRDmamOfyx4TaiOmOUx+xrWZ+xrCscbAfEJupo+pFumP
F/dx5qy4cWIk2T3do6Api4Iv5z/MWU6s4wsvDObVqUHDZcxEA6gFQu4Nenj/k4GmyRGX2Q3/UJhW
zWDvxA6RAkGTq2AqcX+e3O1jZPBU3wBFEAnXvlbeoW3Lv0l2s+8u/2ygWlorf6/+IP8j/bBP3DUu
PS2Ct070PjHHrMxKyWcX4Treg4KSJARsF/b2JM8l/uoD41bqeNkEQQHqZ+hj5Ou2iPhCWcv73S+1
tkVwkCO1H/Ph0MoA4Rne1R2l81vVSM2+CU6/b6gKZ08bEBF/P5bTK7WUS24aCoY4zGWEr3hQVqbQ
iC5+HwO1granNTTTF9nA/6tIZuof/ez450sMkjvFj4HSqVwdeikA2pPKcljmhIDK8NRMSj/UL56W
dMO3ZAwILUqi2VX3GT23bO6UXmcgUs7rOWvGX6ZGuiZyHZKaSEj7L/BwKwt9cSiDJlmV67Y8RtNz
HYxmki4KKqFRtS3FfJDRXbnD0R15VCWwf356WYzxUIFMsZA7dCd4zmv2ezaaw877UaxZ4KX54p8T
GeKL8UZ0rOY9/BnXQGe4YbHDrL3Zz8I3lZt84Za8yCLptYJ8Xh+DPFVoC6Aj4LkomLqM5SVtXxyB
+RuuPDUmXdRv9cjjzwikdnHQ7pHc122OV5ofbqgldDelKzRlgRwV7Z4QfnUwIw88JbSCALUFBDzG
rI3YB3rGhTNJ+hm6lszQHEmoNY4z84aDsDQ2YprS4PAcTKYcbKysaNkgF5v4t+R1QVK86SFSyVXE
WnwrKxfDUVKm9eV+OiEY8bYvBQA0+4VpsOmE3YeuMToA9ouCtfh5JIUajm1UovrZ/4aCkb1fTTtL
qEiMcAe7Ic/M2YYsDFW+Wn1JI6eM0h+eFmzDYa88EdGGPQsYowbHusAJvZdtHJz60Njjxfh2C5YJ
0/lHc3yo832VjkAzvEmazTatJdey09bUIk2cY2P56pMw7gOPAs9KmfB93dNRhdlhRLoDCtmCiMNg
xr7apSLaap6W1FmANLPdKC35obBtMYcTTqlVPQln1KLy6SNcX46vjqaN0DYd+zN1Kyl5XlnGTmQX
7McZkmSk2wux2OlUaUDkWwC9rQUDm8yJBMkhpoQ5IZr59wyTpQgAYRV8kCJ6Xtnxi9If5ua7t2Ef
ROrSvkfI2LmPHRxB9nQAAD9JE2xDxfdJMShA7NIys+ZnuvMn4HJ7Ne18yoDRJ2FBN0hhEDf1R7e8
PaRKgYGLXhgq3bi7yJM2S36f7e/YZE/bJ6mu9dLu31KJU5Kj6kfxaJMJicEHVQZewwnejzxHHVpi
anwRRcqr+gGxHrb3c+Z4UQSsfKZNGNfXptMG4Rmjc6iPN2VLi3vLwQj5LoyhkgCahrhyLziieIpi
vDpNKu1zQmG5FtyXOL9XUaRIBKIxF5ZTtN1uMRMinXdaj3mhU+AtKAes0aGUQYTcpwGXKiozx751
5b9+tdFmibfmryahXQ9SkGBQECWzIblp5grvi9JvRVF0XdaB21Iqcfq/fVy3hmX7OfxbJOjL48DM
+BiQyyzzc8iMNF03xddhEu+f3uNni8x/A/PiK9wbE+ATUNOwDq25/PzQh/g8eiu8sTiiuxz8hZI5
CxXGgSRWu3b2h8auzRlJm6fJ1omEOV59WGDWsQzAvcTbXIh01QWEYrrXG3Pufc9Ubqqcnl+xngW1
EuS/QhGW0QLY0Suo3qxEP4CUcY2+rN5gWklSJ/CtAb+rcEs4IPfIfOsmIh+gs4DtWN3g1owMlMwz
uhaKUhSgQtxDLkKWRx4XdMfODYANV49BJ0/sXgrHgZbd6snNKnh+VX68qdP5of43yX+KGERCFVdY
jCxbkDcw7Hi6z5tV/SENF4SnDRNH1Wl+V6D8cr+WfMQZP6IOrTynfnwMAMgVRi7/fucem0wyDujW
ZDdUdqVXAZv0K4qmPNoylpFIPB95b3sHplzu6nhQBSrF9FgSNbOQQeYBhh2jooFQTQfpi/4KILE+
E7/hbloTJ/21dnGS32UY/U04T/TlcHndZ0DArusaXDKgpB53ejybzpfnEH7rFpmRrJHBqE3LGNp9
3REu1WfD4Eqa93bNO8PxRGfU71/J6khRg9AexYtNUBf8jPY49dwtjR6/d5L16XNMue/BBNyo+r8z
prp10VFglx/VKpbwhP3tye3eV9jvEoNe3zlZhuVZCgYbAkQ+1D7y0FhbNHYrGLpXoQweLZefffeM
osz2bJRfNy0RSeKRTOWAqwoZC3XOuH6Y1aLadkL0qmAO+ZCYrSrbfKfkhZbL7ILm2qSwHfuAvqpX
GYZqRRErD6mVCHVtPKCceru6ExlWsJY06JdtvscdPMtql5N2RoV5dw2M/IwGFxPAXOFIIJKAivtl
lj0aUb29f14csi261dKFLjEFLSNlSMGXCbIhTLh7OnuNocIBVwX4s6slOxUgSLhn/+iH3Mi14Wvw
90wNVBIE+ries8OVilo42A2knjXimZ8WSsZgma8B3T8MhOQ3y538vUjYyNTDTsZcEddODaOQNmVE
AyHjnOw8zYWR5GSdaVe3lZtDOQbuZqBo01H3mtCFTeuIaFhTU7srDuKjvmkOPj2K+5deiQDaCZuO
UGVaWjbNSiegLomMqOU7oTFAqF0p9GF8wE1kv2sKkXq6aEILD1uSmUlsPCDbwGNlYDNC/9W8d/jU
OgRLdEo7A+3gpfrSzuzAgGBo19XOPviOr3sva6rX/JDM4KsqRb5AXf67qfjKzvq6ExB2MFccUuiA
mXMpgsSTeZN78y28dqtFbqe+mjXDvonQNd73NA9EVEmO8QGr/p+PqXqLOwrqHwbSgy7N7908RGBo
IP4yaaDDfJB9R0uTPKqE1IXkOy+8c/BF35VU8YCTn0CKL90D95hKdu+gXG48dJ1NmoNuNTjNqj6v
gdhJtP5yTCnrkeMKTqd5rG+FlkL9IOxjsuq4IE9q/WG+b6BOWGep9GNs28J2D0eoeh3VcQJogJdK
aku0cA+HNb03Nz8fxz6JFUbdFsdHjOj6TPjsW5bO8WuQA7LuGJNZ0+j7aDzEF03Ps30BvRrPoeAN
1cSXJ0mM7agjNn/vK6auWmxbZNYu/FSF+WrKQGpvDqy1ZV/UEdwTdJg2MuTEvETJJcI/16LBR67F
c2nwsIqy6VRKNL4IzYbQoUjN5kNtV1BMotNcHzqGBECOT14d5OGm6CKJT7f7sAhAgriYfHk4oVqK
hLr2dilDcMD/g4OehYoKjNNQqLt6+KB3x0pqwCy3L+Uy6jlH5dhR78VMut5IBnhWmxYYAABhYNnk
JtoYNmPrDR4mHKihjW0hklhc2sNGwFJeHrQJIsxxhF1b5Z/9HEAnhq9xK/SOnZQy/pRzK06PkV7Q
XetsfiO3hiQdxRvdwsEc5kdHwN37cJBYuVVKWuIKVIvZ2zLyaYI67wrRDwMq8FXmOm/r0ANcPDmO
OPYRWdrP4tHzYJ5URVI39Zt1YMpErnuk5grJT0mEHftJdjFF5DIB+viyTkAiZwYrPSDxDkMomoVD
vL8i1RnlroKxgq4S01GPvJLG7i9ZY9OtPj7qqt9lN+oBUxAqnNU3m+oc7tYm/uQUp6vjmZ0Kh4jF
ctA175RCVNtPFcqF+o9QbRVfb+1M3jMbYWcDes8ttpkIKEqJU+fprpMz+u/EHh4H57W75QF6sAJS
lwcfzs3QltHEc2R70tDOO8GoAyo2tR/fe8fDOA2yvgWgch2QLTCF+kR6l9yCkrlrlgiJ360Tm4B3
KFlP5Wxbq97exzggmP21KBvvG97+nD297gYlM5D/GeEKs3fuZWtJm/Lj5EwnxSzRimrNVULNb8Sc
7PE7VmSkdS7GIk4Ex+XDkLt68+6Zwci+5vhHut2bJE3PSmSGkenZdqS/zdmkzoH2S/Q46BKwJNUW
U+5QKP+LT5nbTsrf7/1HN14DngJLGI0on8/V1HTAsTPr8Cp2o8Vu0yjbEMUH+wZHd2ISkDSOG0W3
QnxdA8UMNOa6TYKszQv/iH1j+TMOiAVw8vH/QGxVm7rTEoNdwvDMmg6M6t7I9ZFBYJtRsODN8BG2
OpLoO+8ODmfg2lUArIbPPdRgNKPmINeqt2t6J2+Ooxb/Wq3KI5lZADlBvHpRmqk3XClAGRU9xA27
7ZPfKDMP6ztylWjfxd4vYwk3Z4rKMmYtZ7xh236I+URGvnCt4b6wUt05lNHF9uqJBGFbNmDr5nTd
BptBlpAE/Fp37odbyvqHVQTJ9y+jKhs8VNTsgAAM3m8gSMLBVdWpTv+zVtzLCCPfyHqvWeRYbqD6
hXMRcHfy42ADa0Rw+wMZzkfgVsk7gr/OGuGXEsP0/97crYaV5cuVh4iq8JGttsCWPnKMIAmBhMcK
uWI6q89kDrt/Y1vS4zWzbt93kEsKHELq6SDClW7gbEVA3YCxEPwzQOshuIJLzT2P5OWmJgynHErN
1DDtk9KCniZTE+/0Dph3zDRPbaA0GhyqUAOEHRXY/8UquKvbE/qVsbvqL+nwHSIP+zsy4e/OUJi0
a9QXFZVvpdGplUCmA66OlwqyxdE3eTl69NHXv48+w2uKaUHyLAY5s/sGvPXlN1vAGKFbJzo3adUn
RtLGKrucetMLs2ZHVldV1iAibEGjkplSCQMoYPx6WvBPaBrKZEeLAdmxAAuvqvCCCFUGcQ8cplKv
A5FlHZ0FeX/VBYRE0/w80XyDZVrMjMqP1W2JA7nFtVvd0X2jvAuYmdVXfMbFg0RglmqN5BQqUZPl
3FiDlM+VRVAJXnrQ9Jk+3BsmD6URvUVxmUR+CmBmsXI0z0aUbmUaIwOOnbYluDWpNQOxcuBjmG0j
RegCP4fPydbcZU6o5Apu8/n9IpOmJVKYZ5WOyc+9ZAVYsDahEH/+t5us1AhcepHgb9F8LUPDRmah
N5WRsOAaq8a+mZ12T75pA53+JWNI8eozyZ0QrURQAbHdHnjehxJGUoQtwRA4hyB6bA39tLl3XA0Z
TrgZI5NOO67HXKaBGDnJC92NXJbl3Ks62U0HGbilXNlO0Wq6KqTlmnRtx8gUAD7W541pfW4dVP9+
/l7cIPB9D2zqnDUTcNibSJuk7JLFKtpBpiXOti4HeQeaL0AOM7c5gwJFpwkVjEE+HMBf0CbcNwxp
9vfLhhFC5y4Cit+yoqR0ccpkYIHmO/LkYUUmK+dgMHsXoxMA9hOi9RWX6Wn5AHxs3BFuq9PoLyHV
mcC5QMsswA8YpgvRWwqRmD3TeXSBDOY5lpYPt81MbKcsa4Gs+XcUjpe5myp1tyxmoW5jYwQYAeFt
kURWVZ/CemrOtiOOdx0hNp+Hg/fEMkMN7aIXFEuTldEyPTJkuh1TiER4+lZPy44OUr2kBskRG1hL
Wff+I2PRPg1jmXTi92uXWpMm3FUWaj8qFfh1+jnU5skC7U6FCP5KsYluMF35qYlqur0c1OV50uLr
2hyYmhcoPC9aZ0DJFnwv+fEwGoNvgEahCaIcGeicOqSGaP8sHgEMWbPi1Ng0rubn/SAL8BLTkQid
+rbGf1ya0INcECsTqlAkGcQgKm7HyTvfEkiLpige+SGG/SjxrCD2AClNyGKLTE3kwEKFRh27bK1S
ie5LtAWbWuK8Va2lESqvDnq/Cpg06a9oyFUk+WZp3I+qwXgu7OVYDx1wEZVnOYDsX/9jIMsYtQi4
suX02+yy/B4Fwii4EeuczbPaBvCMvP6XuIRNVTB4xyKr0GjoEkr0KVJhnxG3XtZaaOU4XYfvDl7k
L+idyFqi3SokI9pLJR9t6akXsM+fQddigQy1fDVbMNjKVql2d9QKFRv9nRbW6AR+JxFVzzij0JzS
epF/ZVvCjbERnsj/kcVS+LeUaOo4xYNIfuHl7kmoIcJjftClwNUSmSmru7Gqe/ohQsThi3b60zii
czqQtP/E54P7jVvUGlVM/gWaO4+fLdxOt7uAkEsJ8zUxGUaQ3WRysoaRuBVrBiYn0WEtyYRiHlB9
gl+RhbjzO5NgTE5QGx5bT14GF5kSixY1VvTzhF9gpJaQ/K1FTNr1+PMB+IXbKiWd61wuVSIyXXl0
x05c+huXt8OL8kTbRKtPUrEAWmVMGqnNvib/yGwE7ajUJOryrodp9KVU/D6Uyl7L5cb6Yb2Yxp9B
gyicusRAlUhNavEkmH8zdCoP1l496REUcnQD/TX9c2jz4mu5OWsPdjy3pPF9DIpLOI5aWF9gLZEn
qHyM5VOzVLeaQO8iXjtBGK6hJwzjj0LJogIneFn91cYYkpsLHXIMbEnaGUKTNzJtMBKhtehQxOLX
N5/6QC7XNcVfN0eMfzp4/8AAFtTXMYK6aMrIau+LkxMk8jujzcTfBB0NE8UTW+whdGQZ6CJm3ooW
A9MZMdoYZat/UjJnmrLKt3UuDOO4zsps1ll0GyWVaum085jvjOG5kgPdLFAr5Ab+C3YEdcW4HFm1
yvlp4Nfvx/D7kHF1gE/2r6PRvtp7SztnrAOmrkbJF/VSHafnzelS46I0fFSlSzY5BZHO9gQU3cB+
sp35mOflvz3nLDLJrXHcPiNmL4g08FsjXK1joBLDy2MjzB9bGJhMay3aAx3YEt38DVrYsBq97VwX
5Q2PuK9flKfLUB8GLkzhVcvHhrDZpOugd/sUQ2HreS56PmX0xKmnCKU92tGKZMLOpYTQZAQAlM5m
ISlmytEZ0KJtYsh5GDIfnlN+iPOLRHs2Ld0uSNHZIqLAzyNT8APlzMfZsvpn6GKLRYenWb/nS9VV
RL7U5YLcHuAkhZGTGPeClmeLgGnGRmFpmXCOLlmxRhjwrdII+QMMjpubPHHhsv2Hdqt2bmo1WRhH
Ba3kyh3039gxytviya/yKDxVeNaWpXldE70zjnrVc4Ed52+AhxjI6yjbWkVLoS1ByUShxvdeRt2U
0LyIKptWgZ8i7lhLzCEtg8xIY09Rxbm9vI7ijZjTzQ0cyL5k15laIbZk28+91KG3Bv6709rTtaKU
WpXS/K5aYTPirtCk1Ar9SC0IchXYXmbNWwWy22L02mPoS63vdECXZA9HAGC2Asbh70WzjldLTW0T
Fm99yBdXikMYFKcemP58GHEhh7yvwNLiWgF64g+wl1euoS7zYhXl/BK3y0MVDKhA8qvHK9U/XUap
9vUykFL/mToJRUvdG7IIG1YNhcJfx5clCq9iZcB37hGmg3uGl7MvsdmzVo/xa/yXvJ5dzNcZbw+v
5EKvL5kuKGp2K5KaEUSwXzTCyD5ZBcN/YuCpGMx5IdjG4ltL6wYv8o8t/vpPbL+jZ0Vi5XI5uRPK
UPRPhOmPDJYApRtSDTL6HUTa80dgZL6Q3vsuJVPuC6lJSODAC4vmeHSpw9H22VhD34GB5++8jHWs
ojHVGgxyZP3NoDApiOfHQaXAenJyjyji6ijxe5eCqS4hNqgoSU3fycPhSVciX76yW0P8Bt4pTUMI
1AVHLGjXQU0XXuagho9eNRfH2pjBoJmvgi83n4rZ7gRMAthAJOo2f9rN4gT/HY/dOPQzWj3E7+dN
7CBMdMxdeOhNvRE9/Y+e+wjoZIWZ7/D58aACn8+a7jXgTFfKqffeZNWgWyW0kocbfTyaoE3tj9aF
Y/yA9uygRk3IKGvo/ah977PyEEQxIsZOd2NhTU5S8KrGgwblczQLBSbvT9UhFfbMB23+M8wU450C
D30Y9pSv6EDxAhKpBgjO3csOkkDDsEYNGBq5ojoG8NIMC/ktiYVGoTrhjDuq7sVcchBKbH6+JwaY
cxiwDVjNjVzcSYcsfCKmW5cgPt/KeoVjVqdeqgkKXDolskexOUtXXbo0/L0PKJ8HSbCyse1h0MRt
7hQlb9ao5DgCCIleTm2C/N81irdShxxB1N/6tptdRD6O9UqjdGuY8ybZVckLCwsxwqQqWLqYyQfY
tr/4PHkEWi0mFCjvJWkg+/z6kyzLbyu9trzgsZMpXS/ljZ13YFbt9cGi2rjmeANrYeB2Gbzcvma+
pUD+L24jz7OV1ouFyGw7IM4N95T3hmWTfINsZFFnhf0BQZ7ZfEeP8AAQnCXRbcykh4g6SiE2iZgF
1d5mfAZgFAbqppbcQEnQu3iRzHDZ0tL0ePE7Q1Hg6SOIBD7zo+A7S09GVL7qZDqw+2Rqrdr2iEg3
IWFSTD7TouqWwi9sgJ4StkVEPAfJex99lrkRJqw+f8q7kim147xQsKU+5T6GMubdOclRMjdxM7DQ
mJJVPo04m59TyA+VGvSUh9WJUCsMYyDcKuh5aHephYznI1te8y5rzy/QKmwhI6Q1Bd82JVR9Ec5s
diwLvvO8T7wkIFSK/H6FexQCqZWVFTvIY2QxMO772Na8pb68MMFWslQrwgTAoBg9EqTjM/2POz6r
0vNrCdeQFGoZwcOPnDL2/5hkSp7o3crU/qM8wEFUQToYE6ZNhHH6BK0hge1AoQe204s1WO6N8YWm
tIFYVLrIG+ViFqXWU+OeI8WmEF1c/p67LWrAqXBGwwJgv7E7es8KRM1VcNUHeHPpacefbnNk6pCQ
XUvezBogVDAUKweWUvsGrOB8PPqCHZwFxcxyIRnPXoXvY9Bj+xVAHV+EB3hy6X89isqisQ/K4AU+
dUi+53pYxlkKz3evF0JvqCok9dCpsf3hnw330Uo1kgQZXK9iMn/pt3y35vUokG1yzsVAdslf9ltc
ozcF5j3zmlpYXwD/CzLIbPbw/NOmbaol0oVM5hlGjqqmKij+TG5eM2nJyj1w15MRc3c5Niqohbhy
RjMdwlfK6FMdnuKXPuryddUoauv1GZIL3Xi4ZluRe6WmuCP/mT++7iwD0NzNwHNpTFK4qLOjp8se
c9oFae0E06XplJjXyq+YV+gjCptvq5pWr40OWPcPHQUAoPk6DmwGlNPQbm+GZe4aPqxGXhjN7zpP
leCET2OvOzE4LAHg/xrG2MnB41KUGHEDPYZWoeQHOk+SGNqKuz7ltMuvwoNgIKcn8CjDhSM2/nsl
uNwKs6JmJCDuoDyF9VAA0vo1REXtwSWiXmMTfxM/D9zVk/8YKoRn+2l7Ool3HVvj9HkU3f1kbVME
PcxRCQko5TFotbVsO/UtSrUxsUO19PpNJh+P/l3oSIheNSorKGPqDLQ4s/bgkSX0tJ7LB2WP0OnX
GedSLBuhJ2ZmunbUpLsE7yJqUDKTEKl86e+DtmZmWqjwnYv7fWY1rq0ntSq5Oz2sFDfLt+Ywj6Uk
e5aZSQtWi3NOYiSY0fLy1rtXEzIckKKmYCFXdwWfuLt9z6IJMlzjtbl0tijqe/yBhiTaoB4JiHcI
jvGSeOsCgmjXaH1EcEmbXHSoAq9CJ/oVtK4UQ36tO345lbhRgdxWju6cQDYSbbJ8DtgVF3B+9hkq
IgiVR8+kVg8sUwZWm1yMx+Cet+wnUMAKHrKPE2BhPtMuq6q59EmOWSRs/8wthgBHxmMPdgKAgVmC
rgCuNLjgUWetPdQI5AlhIxwsMP9k/fVY6PgObEsuGlxx3yZw5MrY0TpZ+zIpvuYm41uZ+HbQbNur
9z6Q6ZfWazoypphPMUZzeDLqGxGQ/d9zOs9z69rnoIWtyffN77ikrjiFdrR9FqnSw7BqoOg3LSYu
LyIao7Xh4PQ6DHkxvOWJsvTXM28TUrE6ZkO3of2czuLNXVduX31EUcO517wUWvzc5nzFNPSTeTFD
oXy3OspleFgVNeaAI4hYQMbWfv302oejQZztKE53CPf/4thxFhlYac5Tev7Fk7VESCrGZSvlWwVb
aVQ1BPoqHsBFG92Bs+SXE8jeV2BmKQ0y1zTVil8+yhF8iAaZatZn1a7a+1Ht9zgnR6RackEifBD6
6W0CwuHs4dqUtBT3fzn1XO7v5w42HOZ0xbEA2DCKGw4o5AF7rxrs4ZrxTakervQlbkfRhH7hkbEI
YB6RC56qsyyeW4nRlZjRvzPKKDdvte9PnjvLOXjv2MlX6jsWeb0cyN9XG6/V0IcXIx01Zwk4azui
7TnvI3eJzHD+dw534oVgsSLKu2jLdyr2PRX9wACT3DHmP4b/4bQO90FnGkRD7nbN1FRHOSfag+zA
uvWHRUS7QwXdjeSsGxYSZgkwdTrzzBJJ9NiIfUjVUaklCJsft6RFCDGXVZPLtTXM3Dt6zDBuJsI2
XRIqv/fmtAhUo4kzXEMViB6NMP0gQ2GqhyQHSaNxg1Mt7NbvqccJo28EPsyDmzN6l6PbJhHPbNnQ
X5H35om2P7HXyjmsCh0MXAg519MNThSP4ApoSkYTlJixwMk3rFrl8SSSMDMfH74j9npmtRDV7aue
9vbPdU0dqeGVp/GGHihYoagkr8rA+RV0WeWT06I7tz4rFFCl/H2+uzPZGeCdNZpKMit8/iJTq8M4
34Fw/rL0FP9rIVim2BuBLGScU0lFR4FaoKKQHB4HBV2R7ScHMCVjpPFfZxgQZApLKfqUu0XJsHf6
Liax5mFtH8rwFby9svHjf7NhKCBJ2RFsY7fct6PoxOFNBGGJP5E0gCT58WGDyQUzVi4qHhwy+h0t
cwQroQiumZ3sXP03jLQ8I9zgKSx6J7/bA03ELDhv4/3Gl+BlQ5R7JGYq0qYucxbjOS4MqOWznsHd
uFT74fp+szzrG7Nb66z0N0W1Zr/jTB2icyTGW9LrZXgm2ycJ28WiiZlY42x2MwEcF+iDQmPsyCaF
FeyPwFkhuGSAymEj7/Og5yhHAN48GwbCMDHoDpx6zN5URnrq9mTZlH8QOXxxP0D1wTyX35r/r7es
27z1h8oaBaqR7vZacTEhxE3INVm8RP1Mu/3xnBAa0OCX1XdmgnvyJ7WhR6gRYM3Kn989KSxY9sD2
WZMaMi2xpfPpKrag/dbW3hDc9658TsatUqXCKjNGC4KmDkjvdEaGbw4z8A4ci6GmF0cOyx30OArM
q2MYB3f99E7x56NNnCSn26ucVCH3aaQPdHgBmiIylUfik91qgEvh6UUTKdUHBNMD/UYLKpHkaVfq
6px46jaNel8znqN47OBXsK/1LqVHWJzh9qcWQ1k45atKvEFHTW9qowUZCvTmTOPVAnEhSW5tTwyh
r8+KEUltNubO/6KR9sN1ddWE40IkO6kzKomFFMSWByc7bzGVKk0ZGJaU2W5DhsbheeyoJkmLZkdj
x6lO6fH7vY1WvQ227T+IM5sWQGldzbIJWBMXokjxL1UTkzdVLQHnjEPxMlEO2Kdwxy9C8nNRcfSz
/mmU4XinefQtJ767wlJ3py8j7KJvSsdlxPDwXOq2ft02iKd8SrAzjSkpFzufAL6C0xKlHuRbgBnC
cKVEtIVsTscdNb29w8+LkUR+KDsQc9giPEF8PHwFbaOcNoRHU6nXsN0+214IHxte4CEkzpmD5ZUY
0MH3emeec9+IWPvi4bhUauIkaPNh1XJVte3ziRF/IgJ6OzzCStQXv1N6Mg8kHt9pLHixrf6aPOdS
yOblfO6jlVh69JrUJNR+rS5XN4U9lTw+cHofUKVKTqli5Jo34dedNr/5g22UoSKPEiRD+vCqAlee
HxlZcG/fH3iDv2tPhVnyPk/9Atmx1v9bVAlDykGVo9lGWc799nGVQQNVtcR6ZIiWB80e+dZ/TeEU
H0xQJKKQisUMIEoiYSDhu+uGYUEpu6eD7a2rclT+MANhRbtbFACFMUaC+mcNtPBbr0SqF5nareqj
pcOpeGwI79llVo37RHIzdjtYWQ1OVcJPlXewnrOgY6X/uuLvRFNYfa0fYrKZBuptRhN8cEENGN5t
HOuHSJLdbZy1T76QTl7AM56XmciIqGgZOFGrfRWJA8pnyX+LWDEtR8VVXg5ujNvW3jEZX54+qUjN
6MWSEYXMymA+vGxbCVlMmVMJFYTGUb6vpJUJuNOOrLiUxIC6nXh7x0Z7EdQXHmqwcvwWk5NvyX/6
yZxplfx1AgyD/VBUTGgciOdsp1uDfd207pRhaDe7LYEyCTy1n9uuEo0gp6ClWkIr1rrcBz7ZyMuM
gV+CiPujgyfZyyF6K7IMbhqstwkqke3RBGgjIjXnMLQyE+bTmmlj+wOBOMW9FwM/sbGLlU9Fp1RG
TJoc7vJjCjrN2045p1QkVOsTrOVv+HwfmTJ+aWtSwe6lLTD4PB0Rk/PvW+TNqhwRKOmPIg/kEMZS
jIAbib2RbwS4vKdpaP0Vw5HzvEmtCC9oOWQ5zwHN5Kt1OunO4bXLLcScYYkWWcEA/wR+dckf0V/O
VJ9Xq1pjlxLAhbAnmYZRuKzoeUOtu6M/UVUTPH39juv5lE2JT/uov07UE9C5i7yu+A5uImtkdpf+
Pxd/mXpn9GLdLgsIfmyDqdM72rxcnSRLq+ty7QlBbmsKgCLC9p+ufrbEJh33L7NVIoKjj2qp9szp
VoeLKAt265jGgYAHYq0cR/4WW652Ab8OTLMto4fMlr298Dzfqz87G72rgDHh7GPZJQADRP+6orrT
uOSdZgQIUOGyjRaCk7CMpntwOroH6D/6FN4BGGkovRtHhpxtk4/4GOt5Ssb+xe6p/deV/lVjtgDN
H3Pz+SKwM9KhVhqgs+YQQ5w2xyiGMVHdzynJh63uDRPrNdWNh/MCdlLhvAyMlUo68o0l1lG+FlwT
zye18PHR3dKsbtZ0hdj7FE+IJQSnK+5fgFmwRG2f3tGQl723WvdI50trbOceo/0To2c9CDvHtpJj
bn6ij64tuy9ZeUUMa+xdLuvFBcP09sXCJ7x6IMbw+Qmp1Epcmn/Xq09cNVZTDp27XLftA4aAL1OO
MWjbraperFw60I8EKU9tL3xmhBYTi1qGbUXGI2SFceJIiLoqkdIzMeGeX3lhtEQXjjCFrwYjumqa
sKfNcbgLFc6BCNibh1qvBHywX9EvDbUb3ToiTfnkIbPZv/nKtmRa1FQuy3folP3moNTC4A2Pr+YV
05RKsYH/j7lMGLpZgpgjzNdcrtsTz+B1gxvMSU/AASx/LYZtS9HAnaNNYoFzrBpeMnjLdWyIO9G0
rlKF4ZbszcLRPVb+9YAsigLULG0azYhHbkvcpGS2RoDk6fa119bLt0Mk3bp6paoJn77qTVNVIGon
YamRY2sglsN8b6ZeDObryEu7wJUeHh5pMJckiF+xD3GQEeO1+sGunzB3TqH056wNAhw1ax65aaee
OBZCSqi4R7E8XDlZSpRGS8V1Fgb9ll1lYUuGfxak9N9p5sIgPGdAD0Ouf0OcC4RdMX6xo97DJY9d
oWJLpofd4x97go9UA5X9/rDrXFabL8Y1kXVk144USCeCNfttiWSsiAn8MCCsxkVNZzinBeoA+ofQ
0l57HQOhQh3kKm0iyP9dj3YwPQgpybplyl/QnFNZKdztG6vKBVBHzv7+94g4g0Nbn/h1zvdW2BAx
7DP7KdLpzGLVH69Jd7Xlb7qw9vchPl2D0ymR38ndIAMfBqOMib5rc8pDLPZ0CDgQeUx3UWBmINnO
RwO+QyYp5oBd5h/WtehFVHfYxGTSxzlHkPqgNULu3X7ALoJY8avcMIVFVyA/9S4FwNahpMGRu4pA
50Lw06jjniALgg5PFnsUVgvO8YlVsVHKe4QxEcW2NgYGFlEXx06JUR+vdFImp3wb2n1qxNBD6vNb
a/bbHxOQ+nVJ08zCmQI+l0yf+lNO1OuvtUladIrfNsiYYArBCg+D4t+WeDUvnwGF/NnfvyTKPMqt
h2zKv/XsnC/AHrEp4jzY+t1meEkhvw/pwQCA4BaIpWCcjD3l5rb2TJRmAgNFfq9iVlHwTwqXsqLt
4vSeA+useX4bz1+l+oufP0rWL5CB0qtLO5FT7EgCzDMOskMm4GchFXyNbvcQMMn0bT4JCyB0ozYZ
XSuCFZOCQbrdqVwg2IO8y23W/p7t8hh2daZZXE4voNEHIy2G4PXmm3ENr62MjsMaRZSAnyUttN0M
U0vFrlgpYuyBrB5T6rvXfmoFWo8B0Zwa4T3HgY9u+QpynV8w0sml7KN3ZEQxFWZap3Ni/dMJd3zE
QKsK3fxMwKhPY/Lnl6nO78X1NjsBHdJnGBbnzDpobx+SnPh8/seIfjdASoT1GlBghEy5i4a88+g+
W6E4wyR8nnGtDl2i1Vm4ow0iZICTzLi0GS9eSNv33VbRHMxZtVFDjkyTJRSBHGR/zIbsZbiApex0
qRfzzRzJqfk+iXv6j+FFdZe0P14TnmS2ln0NH1XaFbosIrKLBIMbbfyht8FKvw6ogBLGsJXTRZEh
pWSLie2BD4Dso6ZNpbo1RqpjAyGIcSrnn8yCKBbRV2Q3O/E0z7Kwxu4CkPbWn7/ss85fkBF8v05/
sYsAHAejAU4YaAkBd7JfCgdpL92QLhc4Zy5n2YiiHa8P+axNvW1mH8NhdnzYTPF/+xezHWFKNWmK
BayUAPnrAqT0BY6MoYD8SohRS3XSViceEsiow+IIgTwosQIQZV/+uO1Y+jVO1Hk6hCGGJfFrrdOm
RMOh2HX0luXGBFqqvZZe4BZ65isi8SdmTBaF97LlJxVdAtOH7qCkCH8Dr/5+nVdhD32JSoWyBtpi
Ao451mNT57PqY/kq7nf/JcmWcSliJ4KBtnM1+JINW0gSzQVQ48b/ag9YDK1PEaLmWZF0G6MtV5pb
TxcwkXdHxa2dfdcPeEmb5zkGuR+Av60l6TO9AZ9maBxu5Ze2ntEkJt5Ks2ZWabtXDenjq1tCw5uh
IABj4CfjUqSGRX2vIz4uVXd+xuLc1jjRSbqL4ZGETgqiwt7UV03BiFuBCWIRrnsShYoi/JDit6XB
et0OqyT82KD5/3ibvouoNcqz8XYKBnHzVWwizuBwKAzEA9kFDI3uEUtgWdvVrRdpl7EDNcGFoUgg
rSSKYF9YE8S1zWXLkP63VNxizIGdJ9CkHGX4lhp+01jSHm6YnDPVRCFRmD0G5e5BKGjC56locbNg
CK4meaZpJaeM4CR/t1oh/nrI0+83vNVK4He9F/FCDAq/hNbDL5R/PVnxq0D8No7JZ9O4HoLWUecm
scCRhSL0I9hB3vw65eP5ByI0NSDH+Dv3by1y62odRCcMSJehuIqMTZEhmLMy4cPTVW+CcsF238Wi
q3mQn16snQxEpr47Y37peOAo9NeiKqdJh8NwseqzrohlrtEEmnNrArfFNdYQ4PqFsfoR9BP6sPY2
t7t2eX2RVHzfSkhbbbXw5/23wf2qOMavKzO5TdeOp8zvMKl7In0MgkQb8fmZU531Gjr/cP1aNHBa
PJ387d8+ccY7nf5EribOQ/nLYt+Win6VA8Q49qUOzVcqCQXkjNM9bKkgGoWnQyfJyB45QE2Xf63n
+Dks37tIMHq06mD9eK797JJY37H/nM8+ABtOKcQ54x2H3AnfGUhaAwFkBM258gN0lEzi8WhPGlMB
reNqqKXNU8pp6ProdW/grYkH6fjkhkh0dwKSR6I0Em+EDKcutSWKCiznTLqmURlIRyZeMW/edqIh
6oKl6CeXraC2p55nCDjgjfJA0rQ9c1ME61imJ8QMg7+hJRXy3sYINC3hqTJ34FJ/F8ICcn/fgB7h
YoDZQrVS0SWROsSDq3o170xKccvl4RBGgEA+2+8lar177+zAznFS2agIe83wsRqVcdJ3HIEuQoSo
kLlgjAwax6XE8+xBJH5s7ru8qRM8pv/lhYetKxAT2vQe/R3iaJefcyqLcIXBFWaknCc4kLOIPWiJ
iQOIavYXaRDTWvRUVStAVCgxjVmNH8eITABgc9J2nv0rkNb3qlHaR1XHbOJHBZ+67R6LJFFBG8qW
pfz3+DmzOmt2qhsNnB57rbByWYMuT5fh9fIyNV2g5ypkbOZtcJ1PtQ44xwq0yQh8fIodI6tSSW0x
qYtPxUz/OaT1/gpUMdyCWV8+t1uk04aPBhmCsZekkeyRwp8jKUdkxlrkXvf3EuAp/1dfd92qVjtV
VBuPr57XAUKIJzgyOnrYchbYAqoj8bHaf+ML1oyNRFtOHETR6YwKCLslVkhw6fieps/9LT30vmMA
hfsFQZGfGXcf+02mgAp5F6BfP0poDSYYi0C6DlxOZ/iMjf3xsDa3fOaYMbD/cD9A8kQ14nr7b2lX
0i9MMb6fYGCcSAs+ELMHd2w2s0S1FKDLCxjQxsZyIeQYNDbBH/22xttQG3B5c9CT4+YSg9rYk2Ks
MB/qoERSM5HEdkYfRmKvT2oqEiiY8QHRNZBsrMta8hXFtvBOuLgsCUWVONTFzqlOLYoqf2rEc/2K
lXAILh1c6ATCMJ57zjwL8oBcTkIXOhnrH32PYF9AycERwJhac/7e6xrIVrDOhEneNwRSG2l4BSEJ
Lq0MCgNKO7OwYXdbhqFL/7/wVKde6uW8Hdp7tTFiWudpC0MzzmdKcJ4On2syL4al3IsLFPd5Omst
2uN+BqGSC2jEzWEAy1cKVAkY1YhTkeuwUuohu6dCHZ1uS+1SNoAWlAoSkPFutVZYSPHB4kLmYJmN
EHy24bf++wBKJ2ZGYAYwgDHWrTfJb42XlVcjhQdTgdb9XLdK4+9kRtINiacDoiundKQTL7pBY0T5
GM7U6DZreV7LsxeD7TDElcdHHBx6RTYnHMM5gx/rxfOfHa3nf1S6F8ImZbvg2+hkl7L01rcupfjU
IkmybH8IUeJrmRlBka4bT9U7QJo+ryFybIdlBa95m3dwIaYsWaXxAWS10JBQDrLfN8pszfFH0SsQ
FyfYV/hKKAb/UeDGW8Levcj4OIcfYFOr4WDqDbijc9sNBktG+NlVVjhzKhfV+IEwrvUSI9DbA+Lf
LAiv60m8muOpr9CAuqujMVkQL8KrtPan6p3qzRziJoeI2xi3Fc/dFCVOF3HltHy2JKpow4Mish/K
Hx/NgCMTwF4N+9fa+vlcfVwY+uxAGSruHStmJQk9E2vxZ/r51IACFMvLMVaOCrn5L2NaB324sI/Q
2FN2RR+eDewOTPEuHqr4UfDFxIR21GQT6J5oXPRSbzuCsKv6TeLHlT6RGPiNVhZs8dlYs1rua3xu
lQR0ksAh1hPQsRjeI08ocI3Tg7LZnw6rtWbjZC0Tlc/UaN67fJ5v006/cRR/LofYSOS/rEtCyhyz
CNM/vkKCtSGh5UFhtttn+YmNqvRpMKkVU3c4X382Nqt+HBdl0W5UYGJge9cnrOqs5pHJ45fjpUGX
rrSppJ45akzcc9EkKUrIOqa/o8Y7htQQ9SfREAPpodJjWVCvmSed9RVtFNlFUhx1Q5LqcZ+zOgED
Wl2v2QVTyJ/RyUhLr7fAu2pB5rsIfUhME/YyAxZOwla5+g8UW8WhWMRUz5yJnxo618X79pXXdipx
m2st9KbK2ZpzavTLy5QCXMi803fM+SLlCK6XyZYWYBskPIPY1JeGNCxCrkzsu2Px+kDAF8ChA/cn
UxIAqhtBrjJJoH+Vahc1/jJlNDIHCTDktNV+2lrMqIOyVAm/MljjYAHDRhO2+4+DcPuXr6KorM35
nu22P5/nKROFNFip5rHA1a5i6eDL9MAR1bA7lXEfDhtTXCqn2MmTp/23vW2Gghy9cHQKYVPKP/3z
NnsYIh7puRpR5eQ/IGculvyxY56+sdxZe6eld14NZ2K0TAi+ffRUB+YasYncYZcVN1FzfgzZ6zVE
Q/OItCsGfRAuNfaeiQ2zkGWlo0HhErlthbhE/FwNxQ39ZVMkn/vqRwyqqw3tex5zXrmBiHbu/PCj
aKMhSyACc+GfHTaz9qwaX1a7ip2Ow1UgzAigJuWwSormzkpqB9hWPwwFIOglD283/rBdkkROiG3L
x36IVpU6XVUfgVaoSIVCs5G/Ypc4psyx/fE8bDCkVMoDhqoaonk/M0gligMfCqrgn6eCNOaaS3qr
o8GqJaFsG9uDbRnvHo2HoUadzKeHVIFpIvB01LedKEEkkbMz6ldDviUKzYz3dX/l7wbo/N7YDF8f
Adzg1DQltv2AQWTYMGHxIqR8SHPkLzBm4rg3MY4glp0ZqxA0+YNelteJsXoHZJ5BRDnli1svT4bp
m3v74t6VNg8p1DQBsnmgopos9PcDvwd1jRWkn8PCWQodYsjqsc69e78iwuvKkMYzwcPgBmJMkYM/
jHsdpIEZvx4E69wB68RP5KIk+6PqPMWR0P4yXRqmi0rvgsilIpqwOIayWeRGa0/LHlJL2wfOF5Ot
+BLz/KYa1fo62Jv08mjzGnsFfz3OKVgvSxUCwDCwD5r/TckE6jvAlq/diltAdsHU5gxjuzNLVGE4
CdBDLfc30fOtZScvPQ0ZBItZZ6n/+uGGbWQ/sqfy7pPkgv7ELNRPY9NS97JABOI6zMXR8TukR9YA
rlYCQtNFmUYTKLiYUn4L3DUjIBLtP9tOX/Y4a9g25OwsYjJakRBgIY3jEQBvEG+iUkzNaLi+fLsn
qWCBKc9yV34EOuJA/VhhsTyxwtHlAgw2SpIA4/aoIzDg+kccFTiBQ3tM+CzuUh679GGcTV26/FlQ
RA2vFx6SOh3149Ne7xzCop408xehun33QYQU0D3R8UFR+6hr8AiEgNdrdoppl7A1W9pa9o8jmfbR
/plKXXohEXm/C0rn1nCxtOCqxg43bIH2NAvWfYVA45/gG7HlmKC7FTt4M3GA2lyPxu/MD6Nh2e8u
z0VSKGVnw1lWn9KPYU2H6HFgIK9KbNfNI4oA1BMqcYKnkqVnitxUv6bPB36FYX1+OGaNm3AX17s2
n6lRAOOqpGcjPYfBWZ4ewxmxLhgvlWDtAsM/vyJlF5l9lpkTBSlXCYCPRTPfIqgOLEFnGIaGhWK3
odMtyH5qydw3Cqwtpkctk+WNQJU4DFRrIHKqTBKoY6Jgy7cvtu5W+EVHARavNYUSZ/EnTDhZeW5j
BuzHb5FpM1m5stlvRz+zGloKs1VbbtRuVjgIoPALBoZwaWUY5ldw+5iKucvR+pkogPcQ0mMjGEbr
36NE3R7I0mCi+WZ0eHmadaX7j5HjWmsEqMhEgnJUsORCJkLISD9zSXv7zY3+xNDjIwn1fmyNgqpm
oaJBv2G3OdNSRBuzPGEwpgH9KFQJ884jzIfzYz2P7wP9An1XbVmCTVl/OVt0DPgbV3sZFEp3g8bF
BWa5yOHu+LXOH1PEc3CDhhqG0ENoKv6ypB73EB3PiB1d2hMxqm252THELUkTO/HAXGwjw9KXt2O1
Cxvfaz/vz4fuBfxaDe4yU8kTZltFtyxeVDtkT/V1P7SQHJsBsIzJYmQSvXNUyMnkAFkmHA0TLnS3
P8EVk4/Psl/mF4NqaUFtzXZmz7CY//Nni7pRTJfUslA7XsSK5tetGXr8P9OBxIxH53FzsWMTpGdf
s4oTxtGQZ9XMu8D/JSjZSlMTHjjRyEdOjPGhiheCFK22ZLtlM8z75F9L40Kef6JUIRnI26/1HRr3
1OY3kFEENk0qlzQK4b1R/Xm/LNn33max+JPjhcnDDASQupscHpvFj/dAhTCin6LVRdsjXUL3K8hG
5fBtVbStbSeBemMpzTNCgDWB3ZZ56r4uQ/cLm7wXc3QCBFRDGRG/5nj8Amu+2VnmGP9ZlCaVyzIl
uGX6AFlfDEza/HXtW02lKQijpdEXd2VGfoAy8hj4BPIPQkO9+iD/0RvuTyMzBwt1eHYZmpCRfdZ8
4zGHj9fkBJ8TEISyO+yu2I8ka9JO5ifKGAYtWPMV8eGatM1gVg6PdAhaAz6z5qjNWoE+zWM024Qm
Ha4gt22f+xPXj+zv1kbKgj+hXYWzDu26x1YYbvk8Itwl2se6mV6mIr2dWFwdIQDHVlXEOB8vF3mb
haMMy0jYvsrtZ7J2zKMrM4EQFKLwB/CGVNmOtysTrwX2HUL19oLL2jSAjGaKeUEWQwT9gn2FAM9I
LSxkiiMZL0h4gsgxMETnfVb8NB4DggMwQzkIjp62VPlvumnmcg5/RSxEivrMXzMtIVgm+j9DUByA
2xKynfNcm9TUvnRii/uCkTk9Cxtye4HFRs09mUgsdsssSL8aBw82hFU/z9AYWK/qrf3Dmnvw7OfL
dqWiVZ3wxM3aoFLgUQzqrXlLQllJrB3+HhEMqSBax4orvKkmUCasSynvg9I+TtnD+y7wUgGJ65DI
g5H4Ljr4GXi5YzigF7+iXx9x7UDbG91X29uF6YsLoDGZ7biHAJpeNDWXT5q6jbaJawGuGFgPmPQy
R1uMtPHtqBqEHL+op7bodxDzkEdf350WAKkeYBlQ6vFve1wYx3V+hoZ3moaPYwnPFW7jxLMyNxf0
z4/8aWystV6LfXsfIyiirfCe2XCkwW7gEkcIEt1oRa8oKLMOFBp2IprlW1mxOYufigPPJgOiPkFd
d7ShjQdNtP90RS/HUwc5c8Dk6p1nDsw5in3pwTTBP5yCXKOEkEtlYxDD/GXh7kAysxTMvNueM9sB
qgw4QiZ9Sy0kOeUZsqbYeEL/SXkJByrmsa24y6RO/LUKbToI76XXmolHD7NeLvtB2M3vmdWdhXQx
VfWmp54lbmy9n/b5hikDxiJ34D43kqIA1v1R24xGsZE+G5B0VenQ5Gv9xHM8AYNWAIoBeC2U8jBS
LvrLuCTW4zTl4yA6NuBomE3x2iCjzhP2iVpMmONPvZyKy5vDP+GX3A2LeH9CDty76r4BkKJ9m3GG
3+DLvd+DUkaLlwZxE4c6NIT9TMwHA5rzWpFCAVnUxcZIzVGllmFhRO65xlBCDcEKXf1sKnvVkJVk
1O/g9we1JUBnNOutKZj5Mt0QYrr4nL8TutpyWxErNv5o5hJBZnZT4QJm6FhpHqIJADM+XD9lHLij
IJ5nc3suxBq3sYA7jtZ6lP7rqn+lmYFSnVXhkVoxzjU1RPHbDJngNeQjb3vMTfnw5GThwoyIdMQ4
VTMzv/5L0LojNzCZiX+jJAKOEkUeRxek8rXogKP57CLXjTy/8pSH9dXiqDG4v5E1HVIPdaWBVslt
CfRMDpzMqil/nRVlK75yHgWEOGHq35V1UrTIEiOQt5By8N6bVTcnbTZZJx6c4oK/MBbxbdxnGWmW
tXUU27B60eWQkiI+Nc12TcyOnULaTT1LD0LkLjXhvX1mrI+WGzW4Xv1bZxzzDx1NEvpToMMJJcUA
oB1GLpCqjZ9O34XTGEQj2ypRqUa0XL0kefcgpXhGKlqCgRmbYrP3i95CFdoSWICJuTBPLoy1R6lG
HWATZd23qRZ74MFS/QRyS4hO9oQ0BPqGTLRNir0ypTq86G4gd6ePZIXc1x/0EAKE66imhgvmruER
rvn7Doqnph18/Sej0YEe4r6OAOekQ2DF7DlqPjRp2nGyrASOGdc8jq73E1q+1gvSr9OYjg56d9cg
sfLGMCEkjMNCg7CLQX5bpQHPg4IseyKVA4MEnjoWFE12WjgsIe9d8ONWj5WUrVpXsOyocYKwLCYx
ACR47A3GXShJR5EDEGd01EfQtsIQXEBGNxhxhTqsO6xPGbasYXwQHCDukCKCKVIeP2BXDWPM2Ksn
f2eNjn6zICcfXjZN010acqATbs21k6STZmrw2wbRAHeF9PPwhIw3VfVE2Jwb0c+zMgeRiRy3GO7j
VMnhHep1bEAjZtCqBWPXF0UdvHdXQKw6sM49BGmyaqzF6Mw9WxUEk8Eq8mYNr4hlEnLqaMEHTYVr
tStK1fKHe6wmwclB1wpWBaPGFswFBumiQEaCZMpK084fos3NbekattMKTjLZTGdsMCgAF81pcHqw
WbHEmwmDHIocz+V/H0w8oE31KNart5QBROvhZUmFLR41rm9YJ3VOOmbnBdiYKgKG0d/zrUnWnC7Z
Yg0KRUK2KUwPV5RegcvGvt2jF5QvKDShHoxpeNkt2LHu1xKZwkn38bUAEd/qOFpanE/MrKxhWxdX
kiDMH+XqKC9xe9uKYmEMG5Jl/SGBq/XvBRx2vS2IQYrjhtOPYkjWR0v5zuHOMEwTgVxDXNBsh4FN
Ii8D+M3/tYDBNwbakj/ioHC2pIObAbzQZwmvepwBpHEVOdzyK49MVJhWcxEhrySRhbeAYszAqNEg
PEUzhac4GKjXL4lSWuE/x2b/HhQo7keJUuBocjqZzQvDeZEObi6NwONmmpMR3f3TZpEnQOxXogmi
jKSI4+h6zpMo2WVb5vis0enH7QaDucTZ83JOvt5sBVwN8e6rNL2nBZ/by0MzHwqrWty+GR0qhu0c
9U0HFq89SXPIT3g1d97WY5GOohuLl9leP7XmjH6FNinT+sibv1LNZ+DKeMKXQwuLF5zLlaOuW92D
c46wEt+KvM/HIr/rYipU8whDEwygeGo+/EqWMOMH3RAoVuJZiPXpJ5RYz+tNCmL07XMwwUtUo6Pd
jTkDLJk+jv3hD8k7quHoFd64n+MeIZ0SojsQ+mRRjhBfcO7x6047fV1CCQ5xZ43hP8YmQjrCq+fJ
PZ+zi9EfNomsV3NZLmrb3QX862dSv5BPQAu/F2bIV5CGG7LjBNDBr81VAc/B9ctwBVJj0b91kwrA
RH9Y5N4+uii1aLEBdkEReSLLMNv842AP5rubcnGkcOHw0NxsM8jNuAxy+4TIrUmluL2XKHUymwM+
Pt2Tm7Hbrg2YJnzJnbTaHOVLYZpXgzffCRDLJBH3+0tBJB6x7BmS4XNfK3v38sMxjcVjMEsqSg0q
mtpRgdFc6z5cH/045He12NrV+J0y0FErd5xWH+gTS/YOmhqx9bS2zygaVVguqQPcrSjcyIsa2Bpn
jw9oecMcBHaLpMATwJQtpl4uL4JKKUlL/cencfwrBGd7wDq6TD6wyC0QgZMmlbYRLGtnsUdFMGC1
tGSg6vbKzE6P/SIxGV60PelSdfAdwI5FnxnCMnLAUjVPygu14wN0uO7MInux9OSNG2gmDvhVZG4V
fJuhm7JfYzSsrlYnCpWSOiqyv7TbWSHQB+l4zu1pyAJ/+J7ymI2bSPefIWAFb4I1LZMURjy+oSLR
0tH+cLa74++49majCk6KcntAlqU5GD3/GT+kIGVlpAQNplxNeyCcaaITSI4mQqqmswZW2S0K3rTm
O/lEys5awZQMV85T0rtlkO7qYRnpWRZ8IknSUUeBA4JOM+Q4V2aWqPGTSV2Eb79iv3RtjPV/Q0GD
kJkhsAJzRcwObSX0YTo6hJ+XntYxGK7eZgjccBFQ8V/98Kc+Ldue3cQ2c53lDP0mPrKfFwNLJgwl
nBUvnhIwhLyxekkVXa+AuZDlyuvxEgVaZwJuTjmeHB/3tVEfWSD6fLa51Yy3oWaosBdILBX0vt8W
l/+KsbxEMkfmTAnEQw7ZXU557EG7L6CI3hTI+vWZPy7srlVcHN3VpBK6m7QLtqAMFCtxWlAIPf/F
dFS87x1zOjOevTZNaF2A/pzfDuB3QYiEGjIItVWsVBn9E/Qzkx3pgD2p/UDk77X9OVIxYrO7ntIz
OqEB1T8Tbbr9mUpMb1so2V15wapsK+cGAr59cxQHmOiv7Z525h862nswGH3muMhe7A820Y9QPzfn
b+SQnmk14alDUusA9QRSjhK2mJA5JXAHFH+ZdV7eKhKj4SDPQp0QvBDV87LKZNZ8Tu0dJjWYosWf
U1tJjM8WkuclXsZiHgCOIN3rojsYesbkJj9YrRS2OmSeINOubb1Y8ESTZ9GY6xKtTVps8ZIms0KX
WSksOeen6mN4CiZ8W++qrfPBFJa0c8cN0ZJ0ZmV7mDlF5GAkQidDV0tJ4sxhWcZcPoseFnB34OCJ
7OGImQ8LCdzGLi9VDZhfCTdvmdSXsI94sF6o6x0B6ixSGaQTm8/ba/I/V4RMFekUhoYeGPCa5gc+
oXo8MNrH7Hqrol5GLTUvJh2DUcUT0A1fMY4uAXCQjOwMKNRMB+upL10HI0dZHkueXvKzSTC9oXkX
MgQ2ctiLMQBxmuob/OJk864qlhlcNaXhb1ycgU4R8aVJ4XKpJO3nGUV9OwlYpg7LPEfjHmQwu6Pm
VYXyxLXG4VZzFNYPz0mANopzMD8Awfmc6NBp1P+36FDL7mRD8xxxLSj0iwd47HI8+Kx9jMpsHj99
qZ0Lvg6S/vYIN7fbIcJ9Vpf7t+qjEaQVn7bRxUbpwpHzbLdmcjuU6oicfYHq2e9Y/dzpkVmL3Ged
KP8JmA5JzwhWVu3C6rL+NiqeRo0NWsl0y/BGASuFWzcmlLQODeaAdQuCKnZmAHRKPvJKqKWJM7q6
d1pk+7NnqjCYGmPuHyO/2qKzP1sReSbC1iE2dIsHOlgA1/xP2GmHM4HmxBImbFum3J8grGvRxYkE
XAbXptM8feZhWsPejNJqAA4V4LSB/esjjLoY1QBsad1ddNUGP2YEPgJTXkBdHTAkKsPcLVfTCfb4
/9zis+5Mm3TkeMUMoHvoZuHm7Vvevx/74Dc72k6BNBfEHeL+5a93eI2grIZq40yVHRFE3Uo6NK09
fOqeA3mm4XRbRtmS+LK0kZFIXLv10YpVmqYzJLxEZqBvlSp4sZksPz5AACqwNnPcw7bPAC8jT3dI
k/ABskjrRacOEvrsjCR0VN6Om2yX/WBjQauGfbHbytCnSvXQssP33azPg+PGmKCe6osGoI6qvlKA
6y+yjpdr59NrW3nViz3v16m+XwWiTXpEnc1LTv8mKL4ueFeAX8c1xCjgbxHc1Bi7GhYeVvdYABLB
s6x+UNnjfZUgouu+0Jj+D4SzpLQIy659J7lp2ThsjxlrwhM3ibfZ3L1U5xlen0GCEw+sxrQ1b5wN
HKLNl/uR3E+Osfvrp8BwxG87nW1HqlWYHJxugHDUM2H9Lu1ImqgzEkPkCL3lTTsDzoRF+Q9ayiT8
CSfyScDveV3/8cLGHvqLOuWz+PC0aYqZ0/Gq8K4Eibt3CT+9KrhSQbZgSsxHNFRRFvTEv9cITvR9
OcK4JmQPpFlKXW6FpNraAMSG8k/CQmOiNwnwyAAdj0I2+R8trgUDqtwCOq3UTTmh1sHzjExWVaDn
6OkTuMOTPRTiW/qcX9SgDBYJyg+S0YR5BWGMpu8hKPX+oFBa8Padwn41YKKbRGFKZUk75Ij230gD
iEwZgfzHt257ENNITPPzFdOpI2z8+4uG5947ZjXMJ5+jWZZofHpELSi56CSAFHZ65vdwjqxSjf2y
QzasXw7gyAI7mqe3kb+xnjnp0dOvRrcZJa8F8YaJkgpFB0P8PPrncEWYVNUaKd3LDyLqjCM8T//O
SfISPVN3/9NaniqO7hz/arWuSy4F+Ohto+opHUh/qQy2CixHZH4I5NyBpzY+TFAXCjNTAR8Mspjd
zT5j2bu27aT3Ga1xGE8vybzJR2it3fLBkts9FSIppbH+xrhEjx794lNuAehtqXQHwmIQzdG+if1S
M5TT5oMIVJOCwFzf80Za8XfCaVgwajtvMUCiwIsdp+feoJHrB2vZ3HrGpR3OwL8eD2VcWCNwubyW
FjhqKOTZrJBIMzfdJ9zakCuZSz1lHK78wHvYMaixagLeohLrfAvE9lqi6rrwe/RMLah5xaZ7f4M+
VlB7xJt/eD4z2fegi1FTWmTx5EDIXKT7b19Cqohl3ZRbTSlXSUJrzIagzQLY2VgjTUwVANrVIP9C
AuPHaFC/ducYK+elVhNyoNxouE6KfS/uNrYlvmac2SYiWuAgxot81C45+GYD8NaAkh3NEZYI0hj6
YfVdyY3IbEvAd6iZhnois45c529uetSAMyU9TvRsVHMikdWEFwD6JzyHBqi++mkdge6YDpk3OZHc
njpHG/2J6BbEOlgz9Y60xTDFE/LEToLIb58maKW3YQ1EsQG0UzhwF9y6oZZe38fHq5apuMhJsiZK
67ogM4cuTrLCVp1WPR8m/xLoXRlmegke0kAVK0dA/iTHaiUlCjOl53smsMTMn3tbaxJZEpjVBNSz
ZJLVDLT5xyWwsn597XtiZobem0X1uiZ/1KRLqHaiy9i0WFol4YehbzdOx7e/gy4i6FcYcnX16l3Z
5SVT5bsZEAbPwIWkykXxbW9jp8S+AgFxgDaWR3ks+iWC8+Cj5qj+5vz4XVCMiGa8MHNUmHrdPGXy
kE9Sj4bo+a4a3iGfVjVBIsS3aU731jQcUIDAvUtYuDbxVDrkWbFN0joXUfTl/BeFnRQ7i2pUDChX
1rT0xa8MpVO6y4Ip74LFuc0tkpoejfJsYgm61IC+UUyohZRpDfp0kbwwvH+/zR5I6Kn8UmD0zn5I
LUSXDndqCo0tR/2/zetI2GIkkJDkleb0K+WVHlswh7KrZq22wV0GxMTBst5hGDBDCuXeHXq6RXgL
kC3xemaOy3+vqjgbsMQ9SbmIkzla+pcib+e0Fjt/k/xXqXlSlU9ftGg+J/CJVNaXf1PCBZhPuRM+
8UiSVIpYZoWF5iVYHkdRRPM2juFG3C23DyNldEMlbxckM1byzush5UpVLsgwI3fzjA6dJsRt3SoM
N4nyT0lxx4M+tsjJTUONjEsIE12jwM47u1pNE4bMfaO6CWj7C2E00uCjyGqDxbA40n/RfTVNOewh
+lxbGPOep6PnFX5ocRYQBFQ1XTOLJ0TZ5q471F9Ls3FIjSR+4cehO3cx0X/JlgKfUjjEVV7B1iqN
K1+qp/1bhogKdKXo0wk5OyDZNkUPmHPglOhTs1ARJYDCPVjoOKlfHh5r0MF1PO2Ieed1elKM8e1N
9L9q9wesexOyIMyryIkRscPuxNXbg40/AT3K6m8Sa8g4ja/RqtInDxe8cMC/pYEqyri5cQONsmCd
cVjWg7jy5NhnvK6knf72sPQBWcHRyJ4Tm62t6FeSk5XShFnJzsOoFLyReGRzRrkrlmh2gRwpL/nn
QGX9uCeVmdf6LOUuFC5o3CDqGu0mXsLgvh7KlOk6Dw6xrP4pgFjoliAnP+H02iqEbN8kXwk1K0r4
oBFu14fUz08FyYl7NBP4oMSzROG5C9rIp3GsS40vcHzRKBWiVLJ5MV5CKxE/t/LUMLj+Vfo5kHzQ
3zjlKvrmH0tGWQT8TLHg5UZqoFQ13wnywx3jffkm/wtAQjLhZpizU7IgLnihMq0sWNVrts7hRJ9u
HQfb8xOY1FMhnRqtPLS2O7JH4dVznNwOJnvIOIAIymdhUNhl/oE4yCHb8F/lay7oucO9dQe7Nx3h
6SjnAwN57XMcp803jHZJ/xEvWArfxyQcklFvvqqYWJIer3+V8PocKmF/4q6prZB2G4yznqM0Nq9P
SpQuK46mF8fDOvAgPSWpfJdPSMaFnXjvPc8POn5x3efJXKwXs+z3OblSzQmgi3Yuacd4/O01E0+C
kW8ERKj/k31mN3Dfm+iP7KTkuBHpxAfgGFTz2QnYzps5OMg/uJTTaeisnwxTd0SNGF8tWJnM1eiw
ez9NbmXmXSezK2dXJo4vtVtkoyRwqSMbvipUpvlrXFHaSN4D3H0bN7KR7Uxh6uD3SSJA+Vb74zU1
pR9tEHSJPjh469ZmtAF/A/R3DtSb75PbmXnx2seYFScnM38degcl8q/wyc3gI3ZCW4tsrkLa38BD
5oi4ptyrQ043Q2MQuUya/kXOGSYX+LIoHAiRMGxQ2rtNHgN/x1mZqlgB1bWk7F/cJDAr6gKnomTX
X/ZFZRMCCXoQOxpF3APaNQzON5TWEEUvbQ4X/s4WAfP0vdEL3XlgfW2oocj/lA3sbiIjnzd8V0j8
c2Y+dmgUY8lT1+l1XgaC6WrNVDl0F5evPj/ADiOajS3SYwQcqB5/1e2gwXIqoysOtHrV8o9qKKVn
N2lYw+IRtTMguRsXoYxwmz35HgJ9q1DeUfeMsDWF6IZCftaPfY2BpI/9xxkFyViYllVVyi5JVIVe
unXlFGK7OpKqmQIkUjWAu+It6hRHdCbifN9nVc3++jFk5Hype3b75AOXmmnibEEIEuIx88k05RMd
ACcZzEl05SoAyuQME0MzNOoZfFCTAN0bJDxVqZcLcSI3hjiO0k71SSUrQh1MA8csNk4Vfsezjs37
Ex0ZAOYA0AqCJSuwenxj00+zBXKUEF8EnQu/YWCJC4kOE2Bx7t1/PfSg3+F3dsRsbi9MG+3J9+dp
FbX0Qc2+DQ4Ge2wVzr7ZxkVhWPEgoB7o3092Aj9W2r7LymVdghs36ybsw2cdmd8QdTDzYu5z+F0l
m81TfF84N72XvnsQiAtK3d+40s8HqR6FLAFS8/4YUG/oBkAtNDu9q24ZB1NzDIGHZrYKDpcaTZUY
bgvrRYx9XX5n/PjBESus15289WXkS6SM5+Kiv6ecVJygG9tQPgPMSqh+tsTt1irwncowH6uEUwdm
LMsSEE/pIjIrhXW3u2JbxOwRwBbTTyaUdVsXAzb05Ll06WSakuI/DODeO2TbSPRhGrMxZ3AiutZh
CipUd5b0WN+4S4IpqpWaT4jAOTJt2UdlG4COZiQFkwEcBYAnjDeDMrBYAOvUD8rotlgtHAVcZGXP
N/1/14ZIU0M/Icp2FMOJO+jTgtOOCaUSP8+EocPecNJJH4k48uD7lsDSiHXd7HOJUx8zisFUiLwG
bjqB9kFEalqjbF4aKALZ7uyySbcnEb2cjOmyjRLf6YGz3rOjGka+KI/78B5x9YA2/ZUT8eXmLmEK
JZ1NiRvIqheItxKC4RHgXTQ13KvKRiGHdkYt9DAwNc0DSKBhRmvq0NwKWtHF99Mk03EIUH5va98u
D6vJLif3b0ZPavunn+57g+khsYnN66M6oAKuy8dVgjhrGFnGtc83DzPX6OR45P0/5hW2mel4vn8x
jQ6fVUF0jAhQDnT7NAS+tB6aQjEB8Z+5/wqKqSF2Ojtv8AODjkEi3mWilrTpaFN7wRB+gSfN+F2K
c/k8NznJZ+tGbtELpVdinZgj3y2Pdpiuuhqll5RN6ddVtPNFt485BXMomM3MvBJmApP3wiREnyTI
kcz6E1l4oqmipxG1E9EF+iwrxQekdknyeH3jw/fsCkdTDnm0665vbtraYeh69G5l44onpzjfcAm3
P6CJQ4Fr8iOBaxk5qEUe/glLm7bynKC3jFKZouzXMdzArN+ZihQg2EgLuKEiWjPPB/xqxhhPsCi7
8dJsaOFjolH1DjFe/5UPRelJjj1BzkvQaJOBuSeBC3CRZZVcz11vDD+Me89/ySKKdxoNA3iFjgtZ
NNZc39N1EQmwqnyazezixqfY2KWoHGHBBG79Z3IODuAOaNfrMGAt0FNozf3/vs8V64k5pKQr+lDk
AjwnmoERRZgCYiQEHIh2/zGZkszGAHpjB5HxbMY1yq2hSd0FtuafPWpj4bVCHiZrbqlbM8LNhadK
tdFWX3UCiwNo1HNKMJqWHFUHhdc8JCO6purD7C4dl3Y+E0UoyWjy9q7awbPEiMnDRMz3ntiGAbgV
Rb5+AKFCVZLCa1xPi8/QlwKFoJkH2RrWXghLvDuML2E5sd0Tq8foGQt/OqrKmTCPljq88U7y4SOJ
wUg0otSrxOGjb1aQRvHFDfiFqTEd/yR7LSMdq2m7kshz6hyGrpOmJq4oKqhIFx9B1ARhZB0BzovP
K4QiIzZ95dcMeVFBD4nXYEO+I3zhYFFFw8l3WAl4bfJOBYt9NUR5n0IMmrBiheycuVRdRydF6o1r
3ty+8AqPudnlFJm0VswTyNmzsxixU9iL09aQVpw7ptz7dUgQLg7D456usAyk0Pyydgpkc6QEjAUv
dD7swEEbZGyV3z4q1L4aPXIerhH5HoIqqOvHd3kJmHxaq/cgeYkgt/WkA11rQQ+F1JXPxNUJWFS2
Ih7w4A45N6jjOQ+wt6q8LDZVnUbT8tnkgS92L9ZhMD55MhnV8VGpdKkEjjeN3ONQIQf9e0ioUvvd
5tOpUHZI/rchNexp5/2r55U5oIXRSQLe/V1tj3QyVWExGWaAeaTulWQB+F6OTE6Pc00Oq+V5NZdM
KXej+xMGOqyX2mjRXSHnSzobp1PX43RTMqGLXmal0vzwFeMv46EyFejyo/kBA7ITnEi7+h0Kxvh1
TBA3MBQaZv3rZv3IcT9kDtAfU7Y6eFzOkigk4lNaTNnRPPzGlNf13bnnvV7ywKMc8ZlK48KjRd4H
yxFkwd3kqCZ3wjiUXb++47Z1Z1GmkomRxrJqX4DsNk11FCAy1+gU/Sh8gs3aiDpjO9STj0q8P6Sj
bPlNh/iYPY4ho8rvE8SXoEcwzBC4Mo8ie+dAp7IJ/sUwHVZFFeewaRtjs1tThT7lW8NLLtkX1DJI
sfGO6XRItUKBSM9D0Ke6NkXApglwTfRFkTHAkiX4WJPZENm2MQBq7+BmLF+AYFlePD3EKmQ73hl6
m9TMNPgiHjhdeUa0YyBmzNiAdmrN2qfWurj3BCUT0NkM/qtYgnfJREqjWLNWQJio5tIiQ7Go0VgY
76oaXZVcx3ghB/KdfYoJTf/7sgp6UH0I1QCkERGxFJZrTk7Qz/Zerlk+qnXbQyIrCK1Z66N957E9
gHmbWa8lNCx/CfCNAJtDp/fG275VTwnI0AOnzlFwOYU74SltJHWl9ys7b5gFT72nfUqAR4wey9BT
dCOtEYA0CPjXKobR30BZkaQsjUQnSJ09Eof4Mruc4Bdl8fEC+YISTn4Sy+SFNgdIs/pq1FoySF5o
qMW+dXEv/WyMipcm/C36g9U15Xe9KRruc9yqkycJbYsPH4SVCQkVWyvo8UfXcMDoNPL+szyuYfOh
X8+qfsEsRjTr0VupBBagkl9APgFDHqXV6xXLM3WJsOhdW6HzGIfhzgWuzq8lleZwwhwA59ztLZq2
IyGspzXxLk93YVCGtasfOqJ3KMYCJgDqH7oFTt5ap3+wNzrTayEDR8lyWCqBUzLRCrteLGJB5eDv
1KueKQP48ajljNRD9c34atETIjcGjfDq8KigP39PlWcIA3xG++oAXb5iSVry6dd9niXUajjMthDt
oSNXUOBemY/JYqRLCS5tpkou9ODV1nkaM4FMXB78DuXsLMtBsCWC3QhWV1lTTPlFYO+/bROe11Oh
MykbZL1opLWzRPxccWGLjC4caDVlLG2Y2JVtA0b4CxysFy/Sh1yoSewacOfwiPRynbf5DOm8YLWo
yez3m3W3kuxS3jDTj9d1n9qVoNtpFO2355IZn6Rdz+ULG0//vCTvzisNtC8qOkfqW33BaZ3Che6I
M7s4NHG3Wnk34mxOv9AxKTvWzRMuxaPO8tAJQ9m9n3aYD5OYHEolgcmbztzLgy7efnbFNAp8oV4u
j0lUDX5AJDFlkix/R+SNeUnPsmGiUdjZi5drESdX5X4hIejEi4AIOs1f8GFbW9xj3TuyVxFk6+lC
3H9el8cE0cYelNjF33Kxpm36Sfzp2Oi6dRXc6tGkbXELUnKhdvk5rc5+TI/7Cnqx1efI4bVJL6JT
Xh6UlpMAzBUk2zVuFQMqqDwcsGtOXvBmjavNzhpMJ3WsC61r06DlBq/PUAQuZt5+OR0Ecvzy1zrp
4S/yZdRY+rEdwTgA20ECSM+oS7kgaENlmlyk04kB5tAZWeiLYCejEOkqcNfuMsY2EhX72U9j/el3
yssYvICHamACvEccu9N0N9aHOY98MEdNQlqL+Oc7weNkioRHeG+mlscpuY70mQ43vm7WuVtt2RMO
yWt1/cituATC321bwZK0LyGttFPmQj6v90zrD1INCPPsGwl0HR4GhxguGyczTNRyw52N9zYcIX/t
TJkffQ66PBWSldhZnaQwe8FM1VsXy/9/pzZ65GTVaRRrCKjGob2K5VmMMYGuvYihHcLfpw56li5X
7tAKWyjgPJW15tn7+s/MAB3yaxmnN2q5gK+6dWAdHyomFnm+sRWVgA46Tra6ZeU3JM12cyoO0vpJ
IcHFSvHRVZsGYi8zqFsSchbMPwZZDVLUomv0DdK7XTDMKtENaVr2tHK7Y/1j7o8MUQWB7/A6LTqW
DXm5e+mdlzIi9WTmEbe2hpHOXcVSPAF61xt/LK3OBnTs0kgcEdj/LOsWw1K4o73S7d4eNUs09/f/
it2q2JgLbI8fTCuxTwY1Naycj+LvDupXqDAMZF3sUKhGwZLbxz/Vrvo3jb3dMJSGgtAu6R4HCPJl
nU59dAjpv07W1POJNEZmFso5DRNnjx4cPHX5n7ktQQnjcEcnPwoLC01WjhbyQVr9nc+Hx1lrmwM1
n2f7nV8pSN4ovxsWj9neFbdLF6liMQap3hadl0sJ1Isnkm4WZiNSE5dpt+9/00tcPNM0KeE6DScO
ZFCFulO9zHGO/KXaapJE8UlhPms3Vh0ZebuZoAStaZi38nvqEBk7CTtRshLzEZVNYmGLe9EQXLLU
vC7yve5RN8c3asNYcxOdb9PvE8Clj53iWgdKuncU0UhUtioyRIUcNfNZVUv9u7ubhJFvK7+6bv3z
9kBUlsdAtBNQ97mAA6kpeQcIeZj3ibrrddyYcuo4KbfAMHQf/LIAbvbwHvL9pOqu4Gxh5PBgCMgh
kYWXEPpsv9PMnvShrtFLWNi4aiyLrhdPQ9xM+UR7UzTiIm/DCRTkClDGXnvdPSf3n/ezBlrZpZAl
YVYka5TnXCNxcAjzbnRCZmPBzhc84sqLqzXQ0DS8ll3a3jd0jrv50LNe5gtyTukH5j3HEd86FP0E
oymeeD1wl8GF7KOH/IcthOtscO/smxKd7dPAsw+wxLXV/LtATMtqYGxTq7f1QnKWDcV51LCFM+0o
n5h236aZvszmYojLtWy2WBVB7ctzGBNg/2kwfjwf5L2fwcWQFxmo5eRJ5uBt8R3f+D7r1dgofZJ1
GMcznifzofu53ihpdfIoh8KpgSK7P2Xi4CKhPwADrZgRILwJnuEc5GO8tn0cbUEiZYgNKk5B1u6j
L48g3rEVnHqEwHZks2dp+HS7GsEQylsEwv7vNzauZ6RYvrDFkS+/AcNeXfdO6aD2ppbOAei6Mk2b
m1uXYRC4FpaVLDn1JnBgiW3Xfk3klsWzTCFNc/pGcXf2iFJIOsmz2bbjIBUJ8zkDCLs1Dstwrleb
m4FEA8YN7ZaGlHFzo02A9WQ+C1TBHzTvxv3pT0z3mB4++AtwENzPz0zsUjGAJuhmzNajN0hUMfEk
k6PsJAxrqGQLO7s5tulgpiIxCKuCrwkIOcljyFajQvLwZVf9A6Wpc4izgSZsWZpRg3vJz1Qdf5bv
2xhAmv7/fijPdhyRIEVEgCvkXC/uElmAB+k7enhFWDrnL7msDYNUS4WdGtYhtFlkaTSS6uuuIJzY
7w6sXwgXmPUjn7u59lq448h+UaVTPTrhmCR3VypYR7NY2OZveuV+hu1ZeTOcON9hQgrv/p2uMiza
RPqrwrqbRRaZpIiLx8ycyIsYAP9hG+2C6k1u8X+1FO3RVMV4GqEju9PHoc+sVy0N1GgX4N3AenRq
SIHYMNvlQPt+sm31uhv0IyImbPIGEOQx3Iby7GEp6Jo6pp6pEmwmAK7mASdV+fT7KeQmLoCLoYoD
HCDlA6aAldgMKCl8y6eDvlCKr653jTBmUT1AvI8CxJ/l3j5L9MUVn2RUMr8cj6Ykce2MTTYX7vC1
Lo97VIIMVeklaXGfiG6zluQe5aY/cjvyt4roibraeiE5tg7toMtIyYRO9LTDXl0vjGxOz/EGJ4Xm
A9JGCSSH4pxjdTDpj73QZdjEXZfhKYWZBlvDXkRFjUj4KJm/tPqU2jwhKBbHtg96s4GcrpKyOESw
PSZ2/xG/OZrYhgiDNBoBMaxQLH2dyVMaJAqKDIOutn7dFCzbch3R3brIbtFQErbtVZLNNQJD6Anf
jWt/xM8nfqv5jX9h5/BU0SWFIBZdPFqLwCZB67YWhISxDalbufy/3lTbNzeWiJiwcD6StnsTUyyH
xkMbjt/vOWaYc29eqJe9NRfSDojsdQzurTNWWjva6eJw0FjnYlRVVW1N6Qmml9LjL+f1bjJzResg
lGTz3SUejg6AyhcB/pFOur5Kj9mbszD8u3npx69/Uge3D+yR97BsdOWuDZB1JAUtgjJOcM1umMYP
jJEjCNBtEP+vQgSW9UjGmTUJItd8IQjRChnj4Odia1AMYScsn5kU1jtjNMr14zQHhGftQdfBPPd0
JmjbzQzOaRrRXMjjgibwnhTgdiKz3MNNbg7qWUIVQkuPJLk+U8fILtd2EbFn1LxJN/yvEG6uQbOs
UjMmZdRh1ez/1pYp4yfiKq4WiyzShp7KT16uJJunB2Gw+36r/Z9hTjhe6trEwCqV7riMhvVtx3gR
n2oib5sbvDTPCwaszUD1QMRwYw7CUIaJyv4pcNf58N4aLFDWAzlpgRU6Q12mmcMx7VSr/bNS1Loc
nJIYM90CadMUKnhfCmr20VNEA1pcvd0dTDroIxfPVeZIPxAuPewKgDXk7yqAM26MNmMskbW7EEpl
JGBaIQIGn6hqMfyFXpW65ISYPnipz3Lt5BC0G0yE6EmS23cDH06abmfXApEmnX7LyiBdS7lsZe8j
YBZttXmvsD6Jpbq39B6vWYg2Kb7AINMyA56+VCmFM3OFGGbADI5x2OxAIFS30KAL0bbLBuaqbSMH
urbKd1LXl6B6SfPFLiDPNBBVodLctDyUQqARPwKy2qyuONi9i5N/+V10uPvqudbUYquOb/ofxe5u
m8J8CHjy2zTAUdU0g7k+AU6Ai1JRJ4TzQILaxlvYh1pzzssvyNEmlH4WBUxEfBuMf/ZIaNu+TKcX
lknAfoJHJplLK3IPmjfZTDoxr5rKc8yMpjPyY283tj2Am2rwJIZHgr79P3Zn3sFEhObtcny69HNQ
Gag9LlHjCiGeFBFqiUqdXW/R3W6xfDmrPNyl16y8wQTt6riQ+K97LseV2aAbesfOmZK2uDwlC0+h
iYpxdzY8ISPnrWTVjzvBDc5sJXvbGbf3QJGCbeNffMW8qRJSYOT38+U4t6BPp9j3tvID3+NMXJp4
HyqjkTGVZQ2gkWrcVNFp5oKqSOoyMghjaDBBxFoGmNv6ygnOXXvyvWwbPkTU993hZ2yh1fCYcnvb
k1Z8kPflWD+vFiU+5c+6fDGnFrdjDXDpmyPa96vYIN3uz/eC/DZyz33IA2069phtIlcOcxHXLxAu
9NY/gJ9TcqvacqG7FfUaQ8OGbDU8waUI2JWRYodzv8WwlvczXOJUJMf90YJzwz/DqpeSM29vh5EP
4rQ5O42X4Yb2XVCOepu5+vKffti/bWXn5KDgRsgkhAPCpPfc+waAeg4bPywzi7s9Ij2yTZo7sRHj
VuwoCmJRDHWvWYzxVWULNgiDLe6tI6V8npvBiH181tcUg8wOK33wQevvD1B/SNp00EfQmutnvkVF
4HJP7iMB3GjPXfETgTOupBT81ueiY0gP1f2Sqj8PZwDr7PVba3CQywR0z7Col54cLL0XCugzXaYg
jZIc10PMAEhl3k0HNC9YiTjHJlG2DvkKlIWmx6nl1TCWfZRgc2kpMlR5bJcf5dQGl8EMRu9NGsME
MT8JpWucIBApBSxvC3VDu3z11Mc9SdCcav6vcDO1nbOhzE/2o8NpqBeAw1POnOSByF5c43N7c4mQ
lblosRtDSD/VPSZQKWLWqaMsg1kjx7dY7nlGCa8HJa3Cj07I9st/Ki5q45XxKNL8XSk0/Bwb7QJv
dbRsRDDNtktXAjqtVQXLV7vXYmgYsvMW1XeAOkcOotF9Ahl9eE+Bcbp8t5LXIdJecsHrVuLoH3sH
XDOip7RIHX43zAF6Qwe68bbnptTdxbswZTOwqK8F60eJWsi8KyTxXnZ0raOwMMJ3/QdI3LHl9IMT
iLvIWg+Cp4z6EcugqI2nnjfnkJxcEeYOUbxfDDVCQE/ogNkzg7LpA4ArHoqm0Zi7uJ9AdWD+d/dY
MBx/dZfEnK55AQY8yhP7BZHh3J4tQFwQYBOGjmrpLlNZD0DXDD7btWZA60GPV9NoEkgnhiQTMuFu
XkmnYMOKOW0g9wV9nZFNlTeDYSFP2A6QvHt/87AvNyM+AUtHc7chdklpSQ5ZfzPoqurvinO6S2EZ
gveZGHV708OEn72FYhMoTNdjPWlsZtsTSwV/Yt0fHLlQGW/nZOYAilUU3VDjY+lkc6SE/AcRFtvv
HmymkdB7D38RJQ6ebQ4bCjr6YBv+XA9pXFnhZvA4qOY515i5JCdhDMKwRSNRAd2zMxXWiRbQnmmF
kgi6xEAHs43hV/i9byZ1G5Xbhgux0nkW+Ufju4WmRTpVshRVeDbd7SOIY4LLZZfNYoRpAr3xiUUV
FMvRc47s79oirJYo14gnMy5PRs0OYeUAem4CVRDVrc+MGSEtb+iUQkei5oNF0XGSX4WNKsfo0UTd
WCKbq22Kv6tNoujCIMsA+Z7K4V53fG2YD0o3Cj6pDPjj9GzbJIca821WC2c8jQAw11vc1nlGRrA2
d6jSJ88v94QIDtgosOlVDSkNOkL+/LT+QkDk9AmyAuK3SgBFrYWysUrGgsr6aAxWefAZIFA0Hztt
rTRkwQYqI17fXZZB7+hdFHiBScyNuR2t5g25jmLF3CbmTC0C0q0QEHRkVDuAaYRUhJzwHbEmFSVS
pgPgg+2Olufk7+oFos5k7dqSM5xvO8fxRICBPbyqpG/QBFq9Tgxi79zomRmLhDf0tAlJT7JhPWWv
5/IWcDB7OsRNR5fFHLdeh2wIbjLJVFfHN7Au6lFcL1NUulwXXeULkrRzcEuTjDNXbRsFsz97UfOl
JHnyLwWgIYdypknNh8l3SccXRnLmcTeoSTSUJi0ZWWPeFxtuhRByT9Tg+uamAXmKz0Hdf6a5Tt55
WRJsimrshcDtMuTMm4YlBX1/7bibEDcbC877kq29ZC7Wg9adxlGnv7yCsBV4Yekxn3G2zWIco0TR
9r75DdeI2LisgnpHKDefXzM8GEGEjW4XhoV433i/n4PbpgG/IvDH6Y6FBYyGtwnKcG14xQGMu4vy
VwGwxgHw3a+FlWdGSpSgt3ZxBlecKwZpVtg0oxFMj+s2tzCTMpZfvUyvFBfN2SF/lbLiKkI+DeRp
eYH6zSHN0UIxDtf7s1f9B+V2FqUcW88qe3+Mk0c0GjBq+NqQR0h2cG/wgi5u42JfSE/ER1bGj1ee
6Vy48p+GicEhnEQsjiR0JUm+VmPtOMPeHjrup404KGrGM1xzHMgmW/e7DaPhNqQEvrOCryrED+t6
RhKq9poLPIOUiwwlM9XZBoWhTTE3iRQ2/Me72LsEAEcNd7kIZy2GVkXIBfwe4HqBom+a9eAhM+0l
+2ILBkH7NoXqDC2HtK2OpYWN5T0CmplhzYrjlYIVeeCVBJNNNPJAcMeEv/AZdbOUukeahb0CVmML
w6Cdfle+bI3bYPcidMgDlEm3d8AvLK926YiIhtlndJsCWhBEWLgm1G9gYu7sxY6jTd+gRuZ0D8UF
783E+paEwTcnLxLBnbNe2Xd31GB4Mhb3x+df7E7r+n/hBfs4La6dNT185Wq+fQ599r9J5BOpor3U
OyyJknzLeMVnH/qGHM6UIYE/9zH/1rgT7Ajn+0Bo8W1KRtn4vEMklg6RufzimL+JOF7K2MAmraZg
yN8JNZj1noPZn+214s1EozBLLfq9KDRyhMvrZhE5Uxi6b43ydCEK95dtPcRnWQzxz7P2wcm11OOI
rkkSpqd3O6G84CnS9c1LYm36pEywqvhBhPIRwHfBDNqhAf7oPGYUk2K2qvCFX5BpJGdz/KL3W5fw
3WZE7oxH3oxCTY+v1Rs6Q8b70FTe9Cd3FIE8uGjPDp2DTDZdIJA7nIeviqIhKJgtXRoNbdJpINqT
7hHbVv/r5IN0LH5ks1XhYqCnUdOcdCBpMsvuy/lEvZMlPsL4BkTIURCJx+L3txxAGrKt7uVgfexO
dN28J027QYAgRJGbOzsEPB+CepTRG0wusSGYhjsqPPzH+bvkPCdXbqKZrszef+k4l/8Uslu7Q+Z0
wTfHVlCvKu6zQU7pBxwrmZY2CcS28zdpdo3+5cyCA4yakur1P28ThAmjtJ8u8n4mU3VYKRQ2m6N7
I9tdbgc8MR29G1PI8sO6emYvaatzVLRBnbKdFnTS1RUuLHTCiyjxtJxWeP8U6kKq8zNQDfR8RHzd
JVL/VNNw586N+gb2TFY4tjerXCtiGRHY+De/O0a4TeoMFtLLNLZkO7BpS9wRYMGsQ1QG3dLRUnNv
1tQWnRuppTSIl5ktPeRY7R7thW8QuH6Oi+QgtwvIZa7Yd4WhG86/4yfIryHmc0eRZ1v3wICm5vZ9
55m7FYBYGlK61E9v3duJNu/oOvugAQUU4rgAOdsmyqBxsNWHQbbhvWgaBvp0hmThnqocbwu9EagX
nTeL6xohFdJi8RjuBgtuTaPu91RHNmYmHQPP5cQc+HubHsD6HL6u4T4GUIZBqMmSjPEwXQKW5uDp
A1E2dzO+WgsJ2G1vwtLCeKYCeJwJF5aqWsybxO0NYLGWac7UMe2nL45pVw142IpA/vYL7yXHgdsR
7//yvPAD79Dvjrs5EgFhAOltu9wBywVghsWz/4wdT5oZPZJbm9DcIvtvuuAj2bhUn5JBQdf4J2GE
FtSU3G7LQ2Dcgu9j7I6Pf3MeqrqAl/OCFisZwmHyeeKtOzbG2a3nAfgSHgFj+FG83jaXBMVX5ks5
7bRM8op+idlIrO5LewWmnZupjt7rhRU5R1/DW44dAz0z6ybh7dEwXUMfiDoBJ/xC94XXTQ/2mO0y
CCkDNg7zPehqrCyDlmYx65Ng47doKpVOZSGs3H8XxzT1yfWlSkZEWBSzReXJ/oauLfHuTXccbEwO
4AVzpq1KAyAAWnqE0HFpDSSEUiWqlIz6myXXALwzF2jK04cXkFgMQzgcqWpwg8AXpVslocQBLa+L
/IKGlqNiGM21SEo0Ni0m1MP3R5V16yBvMMc3uB/OEYh/VTOvRCXCrBtJAuC8FoU/vR/9jKowLMSx
4AaV5HMM578iT/zj2dI8kAkBxocmZe/ms56KlHZiNNpOeWKUd975Vsu/fo4cE08CzcXdzBD48T3H
VH35abz5eeTcYWzqXSnOBAfnaU9KogtrTvsdjEGL9XZjpZObK1C68GgSqE9zDti1qnHarvELJlrD
K7FZ+DMbUS4Vwj7nlqBBHy4Q9ZNUrrFzeyF/YKinJ+HV5uKGPrKf3mIXu7A2cusLXKCnnaysSopJ
h7HSwcywl1ZKxKNpVsi6NV3Qk2Ziyi692XWncxvmwrXLSIBcTP4daG2YJa+gisRKXJIYqWRPRab3
rVTQP0Byt2DLYY6az+ejfjzVnOfS7dTQbqVT2ljKB7o7OHP0oqs6AQa5cAIZsTGo/6Pw+EjDTVhV
WXFyzlGTBOwecCr/LMrPPQgF8JICioIbOcqizvaz4Z3G30TUW/K6YJiwhjL92Tp8tbs4MK5QlXn8
tP/8wbBSCcjFVGfLmCihP/B5Jnf78apxBtJ43GSWCdQMcuTflNNiOPNYwsppMcHHhtDhe4DqBMqx
Tv/w5kv6/Xq0gAkl5y5EbYZJRzvIkjISOFyWQZdPWpkSHGGS9jodrELL6G3o3ps3mBeA+reB87fO
zupik51EPUxPHaviV3WHX1fjMuXAlWCd68BDGeC6qZNf0YIDmigDR/zezvBljmZGLUtOiZ29isjF
/WBNjazw1B47AbYxKerab6Wq6KnWFwvl9VAaw1y9XaYKcvRAPqSWpVXUxUjtNrBe8d7LaeDV+sU9
YVxjBmLfbTT9Et+gUCp1h/aRhgxZS6CDaAt3PW5qB4YwmYOXK7Zns6dOXKzq0o26uUb0wmiPm30j
zworfm/e2DxTIhTJDllyUzp51XdJr2KlRM0MKIeJTg9i9fm9M+/gdU7md4lSdT0idyE6XUJgTwjT
v7pBBpYDyAlbwi///Llj/4zucVybnvNxyYp0DCsUQ3YsZnXZFxLhp1QAPVHPIws4ZkcKCGghvL7b
9sCawfVjfJsPMzCMQmuB+0y6NDbKY5LixKdPtpF2IuyqElTc24ln/99Odj8EdDJcD8y2iPDkgb7t
y6k+j1K9R0t826KQ5O/yzh5IJK52ZKCxHZ/CFEoVYkT8836NSCmZbOadfT14x0DhZWoPEKuu8hwo
umx8mJtt5HXC5I/EF6YOm2ssEMCCW2kU7WYJpf5nb8LQYcFHwUNkW76jne/1TeZGYMLs+UuQrm8d
OPl/PeEuXT7+ZLXox8ixOTWDcgDBMEnK3uvAXYG5tZKk3XJoVm/0Tr5npTuyln7WVfyd9lX3QyTh
uWhg9hYiOEhZBhxgHjV6Hy++nT9Ql7q0+29+/1muAzHdnUVCZlPCxP6J2D25KRGCreeZSBzRq9PE
HINufeekblMuLkPoBif9XO4IF0Pv5d7HbQ/rA/fT/yloq8uZ2VuxqD0pjbJOcjdqZ+KlVgn0PJqM
Kza8wv70V1Z0RQvm2zr5oMYIfMzqHukdabZw0L+B+qr3oaZTVaBJJzifPm81ssSREo6FajfkxtB2
hf9WCsy1CEZm1SvMYw7Lq//GMmC76xN1kwk/s9lkKL/Aas2pXSHT91fuQXyRY48+ifJ/N0dHhPWQ
UvjR3OmxJrTkkta2t6TjwOoemf7GwHueBPIdBVD8t3r6eEMB/R5Sl3ovg7jEu1zdXwMk5/EKzVP/
r/M/AYYERV8pMibBFw+M/PqFpP5pQJ5RNRDvcCgh3nJqKKr3IuQ2KxNIQcMoJVIZNQgcczEa4+JQ
ETiDm1wAXHr+qXmb84VpxMbxYLdOCj6048VFtf9xHcZWe039BGHHKcpZMmJbLyLgYTdm5bmO/ri+
4gfktDaLlLw/hqrz9zQoH7H9bwrHzDgVPSzNRtxjSI8QABznzOfaTkEMaF3a7bawH7jPrrM5tnyB
kdDyUo01qmW/m93a8k+nvio+kNgtSj3NKNnnwApbSIVROiefqZz03sfNyMZoOOydTfQRnN72nnu4
vBbx2CCYTPBW51owM+suLZNJUF3hQXOFcvsSxs8E9PxAG/b50TEVQGfk2Vs4xU0OruO+7BX6HU7O
wKw/YEN6yF7W/08nT2w0lJvoCrDtVRHvW9aLZ+TUR8PXtacua0kqkVBnpBZNFLwzQeS16M1f74W1
dAd4MfCUEp33pxxYeae3AssRtYaHr7Iq6fmHo8bMb8phdxUEhc1ut4IATlYiT2uceN4VxVQAeWu4
Y3mLHLTaWAaNH18D5OygrX0TFgTh890VY58CZH8yHTCw+xvdywH4bd3k29ye6+bquPBV55mt7sCR
fanx2DpmkbPaV7AGtvLG37Pq4bJEK35tohY4GJCb45j38BOvnphU0Ry5TwQ+b6UsW8kTQdxD0EcD
Bw9ADar2G0wMzBMDqIrdUzrqbDAJ4KzW1pCpjV9+7k6E8AQrMd3w6mvuL+6rwStz5GvgHkTtvc8E
K9JcN+qRdyWEyQ4r7VFCadDx5/LMbeZxlPSx34cf/LtiYi6imrSacQ2F6YJVsvQ23PmJ7dmEsRVz
Tcf+rfn3Ymaw8o/C1FAXfxGXzb8mywu+X4F/j/px6anbUFd1J+/IBqBm1o3xao8FM8b4z4SKNavA
msWVQS5yG7sHbd30dTsaqTufZusKZ+v01Jv9awNSTS/iFJjr87iQCYHBxqaIfOrEsklvWgv4MR9T
Ei2ZWLxHJ+Jty8ZGeItu/OxnbP88l7DQEQw/zR/gV5BkpYF4/74D69Puy0Av0DZVtI/Uw4qoa82u
BFg5D/xKK+EuRw9NvmVJ46Ii6sVr3aB0oB+btVyVM/ICLHzoJSzCWg4YnJt35t3TcKT+BMV9wMvz
ksN70ilHjv0BSUf9ZXmx9nL7GtE08VaCBeS1Tf8mZb2J7BlaEg3FNAYd43s8x+Mj+OCuvpomosn9
u1bMnAIIJ8Fhk05aBU/oPfNj1RsSrqVjqxWUbascNJyvMsmbMHs9+MaaKl5r3WwfS5WZg5nVezF9
rI33TKhrkvPgyhtrQA/Qq3V/i8lZzIqjZVpxjhEeQBP8Vrqj7nvHcjCHmiKXMu2Pp8ivp6S6IbOJ
86wTEfupJ6kxrOfmg9tfRKln2JmrBfgrgBz/7OscYu5aqT+kGMmexNd4zhvnGEmsr5bf9OVwylx/
X4h1+IVcxhzv5pMaaUGTXEXK6zZ5KuUz4pE5sapY54NeibEvxQFWr9yKlwkXkKQBS2MBbkjSVoE5
LCbP7f1nPy2nRbvO5cLiqt+hZHCPdNpE9TfWokQMjS0CHdaw4b1vMz1BFFFyURc+zMYc2qLmb+c0
5c4jWxhGKgEMhUWdx+d0cYWATR/ucfmc44mRvexkt96o3rW8HcQYniYBBQZE2LBRD7laRpf07/Xq
DT1ln0RPc5Yaom7wN5tSSxWDgCHKt2jqOuIc9SdQfdnLGkTXxkidWYlntzsU0MtnrQISVkUX66Sd
r8Ngy9ifKBPdlEFGTL929rEE1QOL4zVGPgU1C9aboLeHAtnhNnyaABoF49s9nOFuwTkCfTrOxd8c
/ani+ntjK3J9D1sk8LtxhO7Gkg2l4eTyaepltyCQQ3mxXXUwG9cyH8gO4w9LBt/+6oFhGfBl6ABx
KUeItKfFkAyjj7rDnWGKc5g5fqxQYsWYw9kvW85PsXp11vZlr4qWisb9KwOmV7DF6/AM8tMWKdIf
vOFzFCWh3Hu3eLpkhxb13grIcZTzz/+otp4/Qjor79GfVvMYRnQCbSaUoS5dvc4IK1ZolkbrMC8D
grSc4z3lqhjLEYgM16jXp4wy6q1V73VsSMlRXQ/ds71OIN9tBT1HUkmGMmPm2UT55VUb5TrQsGJH
xZzfwOwDplWXlKiRoD19ZQ0R6vVUvbNcdaZQlUbhvASVNkAg/5Q5lJmb46yjw0f6kUpQUBDwOGAU
g19aoGeok2kIekESZ5LVJR68DLwg5Av+uECTYGD8VCpkbtJF7NLLPxYzsurczudhC2C49LUBwOBJ
EOlwwuEIoCcyl0H2L3cQ9gjlgiGDXnli7wiiiBuhXXgz3+skSqMe6O+GfBdU3VL54h9b4MVma6GV
3qJAl0heaYTvmwOSDFLCZBVGRwju6lUYUqTfIwKsoZI7SEEp0mrSXxrn6Nw8qhrFOF6cVuMmCwIz
XHjV8S1Yf19bc+k1794AMdkOG7a8+zKPIk1qnvUrRtLqlVYETAt7M8R73C0OCFfRMjpor8Ibw6SC
bNKsGPPcHzZ4Avi3k+eLh6ILMgyEIvFvgrmc2uuojvuFHdCgivk91vfNlF+YnWnwSMKnbx0uX4o3
3RYmTVGjDmk897Jep9g+XKh33r9ll2NPimyjIUrFNfrzobcg5pGZjPfVm6JOf8PQOg6H2I8AOUvs
uSUVvzIA+kp7E1Ai1avyCoX+KbIl38QwXmojGStawuogrLKcU3/MRXrv81tgV1z7SpTDGoW5055Q
fy6ymdd+t/G3a+s4LzIeebfIy2b0D+Ti0x5MSf38zXj/N5MdLtpcbrGeJkr7E9+zepHKqA8YdakN
hizl67KQfLchLda2qU6vnrdAQ308w/ETUuVJPg+mVNJjLjsFCZCwUuZ6sh30qDAnUSCyLToFylI4
yfhW5AIqulwCHkQE6F9i4uI6buRg50YvZ3OUJDZyPWUBvoXRZGO0ppPuoR3JAuWSvjLorhV622ok
X1/dr2TEwwWDtFelRlsT980CE3wx1Paq16E+gbZJ8fz+i+cAz9B5mOJfheWxNrL5RI2idNcTaV6s
O4zP9337fuuUE6G46yIpDFJ68ZjSlVzNRkC3Vx2uLr7L0o+gPrif3ZLG/M7CVv+xFnHPTxlCeHEM
I9fkn6z2UgoWG8tD2pdgC/DEDoqyBHeuFvFg/vDuCW5tUy0UuX6g4brlG/IzGEeFc2menbhXHd7p
FaHOYwnM/U7kOKxUww0kbEBsZc4+mSX6hgnQV8ZLFUBX+q0IePIfN7oGLmqLa1qyRhNLX+JRYv0/
jnkzgAWHa5FiO3IXRyiPe7fEyW9G4AxDNvS81iOFM3YwPRLI6RlebYjM2ah0SEmyb07uwQ5UgGr4
25DfA9UyRAwS/EQyPqptl0F7fwXEZgvceMRWVKTGXDGY2+Y54XVWaSlJA4STV6shOpDYnNib2GtJ
E3xvhgtWYBpuaf38nHTzMEE3mLyWzS6SybQmPETJrtTnfUG1/NRYiBD3D7yhUMrzO+D4mO/yx+F+
FHK3PndLUYWLvSjdMDsr1UWyzJlQ/gCEW9IdlrzCOKDt9fqn5DO/MPiqZBSw5T9szxcKsOdup2XG
ouysH3gftuwBjA8liYj7qyJKbEWFGwZeMjEeU5Ut1KbzN6xkxB19jie+J4s1oQRal8qPkF1obPYB
/qyr21Qatax1M7pNsIvibTbPMJja4VPcPRrzXC5+k3lszSD/ZyUACa3yvpNZ3N2hCwJAVPLd5ipG
G3lrx/MZu77TnKtfq7CJhjI2UKqJhXYRlMiUsxISEiylRahSFc7MNsRS/csNYp66yRUBixtRS5ed
odIaf7dY61jhEtcsDzcw6JBdhbmro9CnAJlHFqV8+BWAG8XfH7u/DUNl41B1WxxccTmlLunkuSDn
QSzdbHs/bE3ssw3au+ezmPG04od6GV3r8AmPKtBZj9Whb1AWpfc6EDmOG2bEPH8tdAcZJM0NXPR1
tFE04BDjPG7eaE78TJbVaWoKi2m68rC9yR3V2WjU4BrhaV4IR+p+pV8NkXlLne/Kkp5LJHSLrm7m
qT1unjBp9pX+R3eRb+3rY/NsQuyckkRmD2VMBWRAQf98+A30LWuVf/T0et1jaxo2uMyFmciqUII6
9uuBZQDBC5G7/Fd2rwtvThXIxTk24PPmvp2b7DtqdMz4m8cAEmLO3ej7b+lkGTKeTiI6w27jirr3
+h8XpTlCXGRAbd9JCWFHeqgodBkVOg7zwhT0ENjxy7+m4ICASlWrFzmUDYr9GNhS7v7zLonUm/04
wiEIA/nfj1GBuey+UWJcUp3cA+S+9QnhlkqLoe8zeTh6tmAluX3jje4quxYOTiqkvlTTylxvPyUD
Y66/a8U4BG/Y0wJ0dAqOVWLO2/jssw4fz7+Md5j1eO4Gspx4AUI63TyrQKVLVxZpzZ+eyAj4jMkI
AOZmQNt3Ug3ANkdqUhSsYqzwLnqp32OwPeYTJChNyzhYwwB7XWkP+G9J2jLaqJVyWudUF9NQ+AMk
08oWeMw3Si9WynXlFU3V7anH1faLV2IWyYJx60ITxDWWON9ShfQZumGU8nHYq0q257UDnRdsqolo
fSr4bA6adNJF7zq29tbhpcS2PsDsDfbaFxN/3DcH5sxvPCMJBCROLu4XfsqSoDBknlLq20hHEMp4
LJOTjOqKv3UBVGXJQKZlpXUivl+U40KohM+DnQPu4JcbcfVzuarVsP4Vdnc9qhedwTwHlRTzCqLg
NNERWs0BZbP9+UVGTGW23xGP4qtJ8VgDnTHGqwUtP4X1FloTcvp9F0fj54UHlNAR5tYChl0r9h0o
/9pHU/RlNKHwZzV4AkzRYVboeDzQFy3Q2P/xuEZRRZHyt0AkAbtRBmQTJMqJaZlsq9X6vr7wWneV
HuC9ab9LvsuuTpJlZbJdi2RPZ7t4RRQxH9RGiATDkOYIJTcfO9Dd7l2mKUBYN0uG6BIB5yZRHlxW
758xyMp1oddHyZ6ocAQGzHfLduEIZPcj71lmK7rrSHW9ESbQ57P9GFsz4zhwuZgEiqbFCGBhutxg
cD77Z26PSnHnSjErDd0S9dUxM7gYy7g76jUBl6ewUZgyIur2Kqqfa3gmv8yJTJc3UvLwkQwFON6r
xww3dC5xFE0o/FVVEJcoAjkIHbnzvuWM2CL2uIRVfmiT30JHkan8fMwPhjcTNi2DRbs9mCJN1Hk5
lZc/FbLs8oK9y6PB9MTVvKkVUQZ8yEeq3/yeywM8pUXWgb8Oy9ti3Ju7alJEPhUVqDUWP9zKkovd
3UxqHO6yaDDszR5EX01r19w1+rX9H/e3gvlc+OeFlLg3FHXHzJJEs7pWYJGfc+mZU1WTtDgaTPzz
Zb8xfCFdeLugH36w2E/7F1X+5ojl8163i3OSRWXEk1rc8fy0cL+60RpNZgClBY5d5a4SuT4Pa4fs
L5eBX15eWArlyCeu9WAcd/3REP0G0Fri+aeN11o/owZ5hqQj33jMSmNoT3V/XjBY9eE+BdxmbwAS
O5ILXckYrw+yWbS0lAy/tf9BkNdAz+tUhmoLtR/6tOQ4EKqEX8d6Cjs84MCODZZKBL6L4s1geXfA
DVtfOUPGAG6Ozv0FdErRp0/QRGdQPNPus8tUnbxmzyemJmCzI8yCykzGJrim2+rUMGY15kHgjcyb
Ur1joDhy+DNZ7PPiu0PFRfw4XY1bg//mAB8Lsff+QBo+BTs9aR0+H6Q99d0oAtLU9eXm7Bte0N0h
AQxMcld9GyQCy/UocTkG8YXj8hiw1KXEGkRfPAzTRnvDM7vRkZiEwB55Avkbe0O/tl9HpqIRZQTw
o6Ux6D8yEJnkRyzsdNkVlUOX30B+5b0gpV3dqdGMZkPRSokOUWJy37+12h8xmpWm8XpWaAShc0C5
fLkAoPo8Jij+LW0PAzVZDrf4TeOmlgcPnFV3LAfylSfP3fv8ZPNRkPX994e/Fgek6tyFQMmzXNzU
jIzgBzdJSafYvSoiayOlrL3F9OZo/f9D4j+5dchBH/uRp5P+TgIAKXFDhNDLiCfymvLwyI9uoJlx
8lzgWKdqn4YaZNk0rdutS5sy3RZHxfucT9TpVJA1tRC83WbVK0S7iDyybf+Nday8aDGAA7r92WfT
Q6idR5iwoqn8KP/4h+neZMO6faivz7Qd02y2g23scmPCv0XtLyNoi8jwAyHs6UaJZjqINddi+XDF
0m8BMJBHQa8OjE3SPF4zhLNo3qI/c1tANEDzLtr6pf/UrEeCKRz4OISS9/9b4aUMjC3V6h4o836b
6GZENTQbbutjZrqDeZMRSqbsJn+CXfnoYu13T+oS5maZsWZ1flsOjhYkCbuPG7R5wf+K3wSK0cal
VrlCBdRuortVid2rM9BLvvZQ2ZuaGlSNI5KYPZ6np++6i2KixxTVlH4hTuDrL9lb5/JRWEE31AF7
jOHubx4WhKCbRvSaMYEToscj0rSAE1Mz6rPj9J6U7malxjQfbh6via8FWIWPB32bH7Gf8AZ4H3Iw
KBHvK+Nt5MdH7THexGbZ8AlggQnK6UQvmQXpNiDWei+U2VBMAaYjDOHKDi/+q1mivwDml1Aj4GdF
2cd3eif5AtbNwlfBN2RZnJhqma/ytHN6K02iKeiI1+dd7C+csDW2uyPaZIzvc9Y1EAnjdyCzwffZ
t8uepCd2dWXsFu12EoROfZnVmsnLAXTuuNDur5lR6q/PqAFperqK8XI0TeQPzZOaU/+Fuf54XnEx
+y7jjaRcEkPZwbL1eyVVkcYy7c7QKnMpjBfPrkigpMSMTRpdGepC69FHr3a86uqZX4MVJ5zhbMgX
UaE+Z54UrHuUXDzNgrKk/hwkk7TJfXNDyI87gzI/UfRTG773Oj9rxHmf5+3cFNd1R+54A53tJmwV
sXTCgGtps0dMaJ/7on//JUvIRuXZ7IxOMEUJpPi6LivKVpll/gM1eJKJXHXOlcCpPYC8ujEBueHA
NAL+gcToabB2dWShmzN5TeQ6Acx2gvGkIuMl5WyEbSTBwvHBVEEeLS15x+Lw9UE2R3hi4rxXwE4m
cksSEluNwutEpc/anV0VY7wRu+Z7lam0jlJC+RzcOtWTwjhTq2BdnrL0Lz7tN9RqyoB+GTKph5IB
iCdwAVJNG+GwkPI7Hj79ceSQX6QoBsrHVDkjY2YWB97KT5np4tMhro7dTEj3dCKyWLcHJkxxZ+mc
TwDONQYdl4AQI7SLOCU9pqyht2gb14knr9AGEtnxXVzZgPlCIY7CI+2KHQJqoZ+NtR11qpRQyoRg
uuSOsiltGKrHIpQ/ZO2pFoiRrYlZyZYPM3IYOw5pagvdrjEuNd+KRr9FfMiVmP2augiqLlhJWrRJ
1xNyFa7wZ3LNsMU9VfKnULyxiIML8oAohNu/IYWIjZAASl23kUgLYGQzYTFXJAq75XzR0EsRKpN3
1MB3yLzF7S63/ws0kSGepekwjlsXZowaN+g7Y7VgDWSBt6iB72xdtRLqrKK8Ce5H8hMvFMJUn8m/
q1qF8NbZid9oG7o0n3HrGkintVNnm7lBncf2hKthOQ1Ae/JM5MLqvJFysuMoUr9x4cYss1Ph9KeL
cPaedAMXWfedrwH1dvWJSJuhw7VqdmtFN3goCJkcA5d34bdU3xU0fAbncvWAFHKFIuCaz58ll97x
Ur1ESc5H9aXMsPs/tAHsfy4vbLRABCNdVmKgo2WyUlVMVz/sdFzW4Nyi2QarNfI8U4a5/pyFZgQc
NYbRxebAnB0/Wzur/PPaJZdaHilAiEPoxLDG5cc/PcwNntwCQB6dcG2fZ9gylZK1wEADoJNlBL7Z
ozUOWgvO25MbslAxYhI2ilxsGvVfIiTL0AYdp2xiQ4NFfK4UoKX0gsrgteJgXIone/ssz63rkpQh
xEbNTtY1voREBaGOSsT17xPk95rZ8omfx7oQvqsrygU4CXoclwYK7OE/idaXDelylGP6cE/DxFFj
A4P6+bQSOFzY14Ux0kEyuYNkJkAZXA4jAA/NtrnOWgEb0cEC/sW+Mhpv/atgsJzT0hvbbD/VVvPs
BnSK4xy+Ea2R3sq6mBi3ml4mcoxx6hmg/l/+zCSwhuTrnXGGNWmFC9+a12xJVHwJnQrOMDP87kSl
kyP8Sa115otLETuNu0EqrIAwq7eEO/m8oTJEco9OO0LrsGhjrhcwbD+qe213tt4BqkWZFZWT+luY
hXAvsNZ/Q49NXMRE+qsBwnGrORZCAdbqMLvf+RIEb7+86toaLCNBrxnfL3RrjN2RQDQ8dstVdSEB
EjPxY+9A1ito48dja7P8UVilR/Ul3xu2Lq+qqILhgzkBUkJNZhY+NLr/P7mYmTxHgc6DMMbSchBs
FJq5Gz0a4J0kenADpPW/AfYOXMJedbIUXRkQ0+NnU37sFHcOrj6EZ1pIQlMIfrBQ3RI7lB2ChPQl
qDjkPHodkzbt7eI23s1ViwCILbOn/2d3NLzSHYyW9N7JhUrgWtF6k33HH2rp9botPMVtnlHMqao7
i1M29gyWp8FN2PSilrGwYVLie5CuxjBDCLg2BPXfltlcXo4oNWWk7qCpf1HOjIrYoi36OA1XumUC
0fv5p2RcRO5s41h25dMJYYF5HADiY/JKTDLSEoUE34SOUrQ4IYebmQgk3H+G0oytFD5CZ/80PmBa
JrKGY5daTRDIGpvcyVChZOOrnxJ3EngLfRnclnDjK17ll56GPCCFwuCcY9K4cG4vJH97PD5w1+1i
PIigty7zi2HQijOD7t8mhFbCczvsKYnQVwBMTjaXV11hrRJwXTP1gCXTxjzS25eQJjWxm2IuWNWH
ZAuez75KuDjvYKIVaeXCsqlvco8JCLa0v7LqggZE2wWVgZdTsCzU3fOfx8ovQywLDGQlaUKKTmIF
1UHBxKBaqTpLoUpOURsoPsU0wKIiHtKHTUBp2Oc8Z7If7gA0yDhuDQEYSJEROJ2jUq31QEGTs3Za
KnBF9QpP5+PqcZI3huoZbn7c6ARp6RA5sFJVohQSJWpQ1DsQx936Kg65x8hQcklz/HFO9H+dp+Qz
YJBUowKerfs/KTRuJijhPiAbkQ8g82rwbQvOrY9kZsZ0T/yQGeBdnlUpi7rvaWijZZkUxGb8C+j6
rCg7y8UryqZms6ywtJ4a3cf3f9MuvsO7OV7g5btS7BhaaAnzNm5SBPmifEg2Or/R7dSmNNJNb5ef
esEMvkd0qzGJo//8EBv/SrG9mANwgHabmNs0BocGl8f/ZRtVwJyLCpD9/FWlGqYVkaVMPn2gV6xU
9WzOflJ9y7rpj46N3TzrbByhAXoRrM1gI+5+Bp7kHfIwIUR2huHzrNaDUoKW32h/hllZO2MbM7zB
XVlJS5IcPic8UQAqM2sBRSYvTgigEH+FOsw9mXnemkH63KcCNMtRUyKfYbW3QLHF4QF+Vpw24U2k
chgXAAnlF5OjJH++Aj0aPeI+ikQ4LhrGr7Y7in6HMeoaGChIWgPwlikt6ImaCGK3/l7klwPmXGRE
HZJBPMhyYoN0GIFzEnkohh8Hzh1+oJvCP9eUb64NRh05Ngz0OxiXGCigkttkRXoYeBCShXJOIg7c
bUpC9kUacd4+//4evrXbajNrkDroQ28EJJCbus513z6AQUefoixSj9LMwQTUykX+BNh8Q5qHOfvk
zTzFukYr4Ft1c8tgdNkJ7UIdhO/9SWB+EP4G0cATfBMGuUkcB9ZVexRECBBWpb1jThG8DZxuN7HT
2DW/e+xJAC9Fa9JR7PYaxGdRliSD35NZUhlVfToLqTbH/EokHcy58SqCsjKfvIfMdy8uvuQoio4S
YDqli7Y1qU6tAsb+knItwUd4rUMtUKmAAjn1EEVZBMrT8sHHtMkz1HISrEiId/icUIzcE1Oq9O2A
xw+c291da+K8S1uum5+9iLoRWYDmosK8vOW6uIWUXd+pQat1ktUmZJRQmFNdeA1n/lho8PcvFY18
JJDdh94XNT4EsoWRQxgFuIZA8LapIdc2dyXamMk7TdACwwy3Kz4H5nZfuwlDshZK4E0fIG3SUCPT
o3LHZTd+PiYoKOmp/6JSBn+0Yj0moOP4K9t4gVvYuoML9de+Q7xOuEZ6hXE76KCuyyxwvOy8aIc5
96QAz5kylwGCtt/iczb8KigyK0rY8Vh9LA/Lh3ybk8N6UvX/8HnyXqJ6+Ex5qcjxU7ujwRT98G4L
Xxgi3+f6EBTvMqzw004fs80VddtQSesWpeq6EfCHGR+SVnL3e7wqmyN6ngQ/sd+bDJlfBxRzOYQT
OaAdguUge0qKzuDBgv6RmhgZEGtHysJhi0Uxt46LEirDQd+zgsQVxJ7vBTPRku5SHLOjKuEtjhJL
t739vO0F35jCSNBRpp6bLra/qnffH/xU+HnpIxgUV4uunfLX5qpyHm6ZSd/g4us/4++G5vPwGnuQ
Ex5P5u5A4u4hVXS0z6gvxM/9sJImfN61gaPqgI/BWPyTbYvMTiq3w7q36R7ylbVXqsPdkxAiQePz
rgRGY5LxvMG5QSg/N9gnkeZqlydBrv+Y0zgVyM5ST+vAfz3m+6VrIPRe95SAFyrN9d/SC9un17kW
Hh19q8b4VysTp/duGCYjQ9+Wj9FplDfdH+We0AW7wOOWf1OLxLWblFxN5EvCK+yT7kxViUoNJujD
vp/gCTH7tJdRVuhxKdlrDjkOGu490LzUUTkvEjFpTOa/5C9AIClnU3eILxYY2yOjyNlQp7SwMb2C
966BKY8uCAWqnMG0b8oWkWcraYvMBUpbFI5aI6UNjA8q4EwGXo/gvB0IF0ZVZrYqcBe65XmmSZlz
5WXsjdXMdI/KgB/nWla9GbnKblvzaioQYQaoszb+WeYiqoCm9K6A20netzCLH9qSAEYItyalT+W/
cistrzE5Z5nDmoq8h0p1bgTC2B2GGNVDEc9P3H2pzLjpL4vUBDjfXUEoTU79a6wDP1bHWHPXmj/X
0UOmXZ4lBHX3vLqSwIr1lUnfd2tfpMQVGKqeH4BKqN02E9/yd+V/ejD7tGFUnVXPRpoQZI3zDh2H
V9/WYAVHt10c7uxT25TE8z7z+ynBCpjVhdbLxak9JwtntoNgoPPdLNrGR9ELR0vqfg4cHucu7Sai
xb0RSdvGkGJAPh3Ww75zM0XEfKUtFMa3fq1gDYK/ktSEUxbB07ObvUHry4EfILSo9FfmkR3p4wbP
rpyi/qoe+RGr2uoXFVe31DVWYBq4NB/LkUAkMoQ2wqwkI5YOqMArmb1aAvQ5spgm16CHlB4/GTqv
U64HyVL907sQbYxus9VHCnY1XpIwGSRYuQQjBNFx/eIpiY8l9Wk2IkYhfgNZN/nqJNDxTIXRLmmU
8q900tD+WA91jqQU3ieJHG9w6HTaVeK/oxvixATLwysdi7d3dzmqIjQ8+qsS+cQafxpPAzCkB/Eb
BN7SclquadR82CxbkXCxobGy4+3dkLf4Rz/3eWk4Db0xmK4UlgM6fSJwqDT4a1N5hI+zs52LRIn1
AVSuM4lm1wypIkYw8K5IXWdrhSUq8VdrBCc649sqw3wPZRVVb6Eh2heqhtW2jzgtmtqD8JXEwsXr
sazDG6T15n/fAIAfiBh6JxwmFqRXamAAOg8OEGHRkAgtxFGdysJQD9iS3gNUKSbNJWczQKVy+pA+
HE5M4kzWcKQ5yF5fZKEh7gh3vvi0ZBwc6BaVxH6tlu7FamFh5iTwDX2bLIuL3C2jH949R3bz18NC
t9IMF9gu3JNSAXP0d0MHlODZf9R1lw3bUavAjs7yUNYSC48kKXOSs/qA9GPYbhOeyibKTd0azkr5
xb+cNcs77iamKNXWshiMfawJ3nDpeDeZaxDQjTa+oXItpV//daRw83LMoR2ShClG1GOy7byge90O
fgTvHmDGpY/TohqcZFm+gqZ28QH4Av6cyeEVnoEg+NlNWR3FZBHrqVbmwqxlgeOdU8gwKeU5SxxM
85pg4fniBB2+FMSz+Gt2UIa1lqkiZ2SmZqCRjsG+5r2qz2seRG13UL4umqctVNlksX+Mzxt4flAs
uKMfWJhS4jPP3zKWNNOmPbEDxONOiHQxOX2QBI6476qP3R+oIPBr6n0iKC6usknAyiUC7QELJL21
G+4G+W4BuFCk8jr2iKJvq9c+7F4ZrHe5Z3Vq1ndPn+PnCCTxPe/Nx7tv/Qa5eZpacRG43sm+u1E3
rtmCzXsPV1BXmajg0Z7O5+DTQTsypY/cosu1EsWt6ra2N3Jrt0Da7i33HLC99WyuvyDuU7p4dsjC
cfh69v2Uz0L6IsY9v6hjO0InY0oaHqZT84XhYTMsyOjdErgEw9QW5F9HesCjO1SiE/x66nW8hmaI
dxlbUYbuAe+ENhzXyiJiMVDC3JljRTVA3XotutSe9G0UmuiakDoRGci6CXMmLzWGPzvmwFUkTaUV
H3d6Hm31fy2xq2vSEVfld6x7KIbQEYFt5fCq6Q8LdDcE1iE46J4ugmKJhpZ6q9uk2iB8KQaZUepu
B+mjBZhwXKK3Hoq17LdrD3EYii/mMw3NjpEJrKxkE166mMMUvyH7hKpcPcu21DP5IDXMAdNTazkv
Jlcw9Id23gox1omcdUOiHEV+0XaCPXcVJT9bNmrTPWEXBtvg6y+xxgHtY9N4JOxAZdNRvsxYzXE8
H8/hRnvhVwJwwPped1/cjvCFQouhTR4o/UwKL4Gr6wEJoZK+J5ydWI3mMxoH+b4Jf44cNXXRDMDk
924tpacHpIpQc52hzJlJmb3VouPhoNfaKO1+a7XdUc0P3N1EQX21QeCGl+lKtQtHatzMjkts73++
2d2moh6cV0F+5cDJ49toAhhsx56ezLvMTT6fF2GL5dnbDbm+Du1h+iq3/uGuD7/rbsbPILfx14AA
3zHkTWhBKmQEWUSeyipno5wUjSmpps84gpqYB4EVpQwo5XwUUEtqaCxG51aafa7gTHIhU07E2GOV
bZhi2LPRVnfyQeP7dIbZRFh2/qR/v5g6mDJ0oOUoQC6CnuE7glIgPp0/2CT8lkGRzv8D8NP20vnd
dFwK5q3xP2QHjPrMTz7Jz+VDF3IkvB53sLYZNRH6cTDg+abakGOw+6goK3FGfO8AxEv4rXs18inU
/ceH7V0fKGH46ebVJowvlqYguH3TqcuwZGbGc8DT3cYQygW2IugC5kjUcxHUJqL8xiRhMnIV6wJs
NjB/zUd6FQDi0mgT7hUhcD+lhicdiDHZb1lDPM/aO+YRYjYZpAQGVUiumYwN1KurwRPfqIBKe6+s
HWxET/WiDCxSReAdqnutoNUYE6kHrrhVIieNeOZOR5SLKRoQPibeIrT+Ww+oyce+Updlaxdy7kjx
z7QMqB5J4CyJ820pGI13MMU93ZnNNbRW5ZslwdWRpG1xWApblkoS2krHHZKkBMMdH8hJnotDbD8Y
obR0ad/TwLKiBzus/jX4mBL4ImSXUup2I/a+06LmlvtpJq8+Vh8CgXgCfX4a36Q72ODhNj77tGA/
O5H0VOn4tLnn57rGjXgyo5eqTC09japfIkgT0SkCXFDvmvOAF6KTHd+gNod9WopC9NRIB9ZIly6K
cgrrV8ExArpazKG832WDhI1viaM63IfBP5URDbB4wYIuYP/YxNbZSr8vxuvxZFmIDA2vkaesrSZt
6fD7Etx1O0JCEUt4M2LIZ1SmZH7XiY/O4IP8cZB9j8AVR/Y5XJolkD+2kfTouISfnLG0bGq3M6xZ
iZCsPr5P7lJ3j/OxTeKQuI6P6iOsD6MTJiKqiz0vipL5n/0WXlMF8CrRPuYoHGHnOKawVObjZQlR
ljHUmz/R35XTBm6YM19nUnzqy+QDcy/6vxkDIaZBP0LV8y1r5Q9AA5rkafjRiG1FJ2bQ7guDaPOu
lYphu3B1AswW/AXIs+0epqNJBVMLzbKISbsN1qRYSK0WTaeeusqTSSLpvl/yoTDdedNUlKBz59nj
+jxwv0WRNSlY+nY1kxJ8Dk8d4m76rHhbK96SOsx548jcOkhi7YmeLPFe6X+PZEi0Ak0m2Gg9MNeB
vV0n+mfM8Z8L18oK2kvJlcCgLH6m7Qydc71FZCpnZ4SH7Xn9QJpeF4ja6GucWVi1Hxyx1qUtu2+s
qsYiwZD2xrifKMHh1tLKFjYeDdHoMoslg5FiaDlzK7Vae2zkwGTLUu/MNXNHYjEnOdavnYiv6oJ3
gMAH8XpGdyQQ3lkzOaIU4ckPoRglqvon4kIieTLO8/JA5KlQK/FCiUr+7YoJM5s5p/Pi3VYSaCyW
lYA9EP+HqoOFOWhUFsffEGSPzGsM9zfIqLNAxpj5uqTV3a7kHqcehS8uqVInFL0sRT2GqX/tG5mr
SvDC+s+7WEUci4eMCTNUvTXFoqgJ1UExPdO5xI8kgDLBlSV0Vb1QzW1kFBIdYQTeNkedHzZ13hIm
HhTlQS+tdnb8prU3I0Bcy/Mg9eiQF16XwVlb31fBJYX8qs+FO524RHUYGWAqHDB1P9ZamI2qROsI
8uTRfX7Ks3WFtiBqxuoNylkknID9wNOfe9MtDRVdA2FGyKuat5MQu8IjU2LiVe1vsSrnlCzCiGgN
LkHXOrik3t/R2o9Q9WnPkJcoAVcMzpSnON204BXMW3soEATcyG5n4h2yg/PJwWq/WZl7VSIEpw+Z
UKdhpcARan/QwpxIZoHx/TfMHOaJxmYOeQ19f3h134MYG2w/MwjRjeOAJa/P4FGpIvmCxWS2ABmG
8Wg5X0ODTDpN9ti4CXwjUGqiggfN6WT1XlqEty/b8Pw7yk9afpsV+c8ztQ5Hb1KqgP41iA5gweFw
/uXI8yAReHECSPN9T2iUr4sys57vlLysISx3Glr8tPC8Ch+B9isnliVzIplJSdL4rpvPXbCTFyTi
JCdwC7KjlDjI4fz1bmFO9tv9TaDlH9d/gvxMOVxrc73tYMkrjaP3Q2K78f/qC0P3+C9LhtDbHPlB
TGzBs6Yem0yjwcFGSw1TaKpxHUNWxkorXflUelZJ8oAHI8Yi5/4NzymMXXrz2JtXbu2geeEIuQ9R
JMJcnh0IgVaKsJAyCeqYAxLx3qVUjUBbGudrJ88CTyE6WYFxlPnFst0WSasWNvz0oCOJA9quT/PW
B1t6tfbAgpjHaiq6gLJ9CFqVvkDIYXNE+vvb51rthZ8PjU5fxYZvGGH3g0Xul4zkOgqMcC8ugRU7
WAbY2tBJq+777dpupC3L6YLp2n9de9m81MkkhQVYOGEIM26hnCTBRtgQpqaZVXyKTpyMDPpNhpVG
u08aK1+E5AbLga9VpGl2A00OBPlq550cTLdaEVRey3GbxS0JShFJCyFWdNG4ElCj4RY4uEnLHYsP
qzGlRyC3NtwGFRr3dHbHulR2V5bbwJZrpgeLp0k4va3ZFkgHLWRKeVvPBMo5tjZDjqndju3upwGB
YngKwsKesbOcuPx0hvbw1GanuPKi8bYnSC5ANRPi8TLUUgzS2TjctsRYZr3C+zGA9rd0jO9NERCk
ulbgTVHvZz0PgEr0bja9P8SQ0/w4NBe68PAum/2rJ7VVy49heIOS6RdPC8t0UagReK0dtMBb9sgM
9E0eYazRcavCOKckYUuxzy6HWtEDVxgOj/4j95qGZ8O7zrloTGur0KyrYctvso5twTtS71g2G/VH
usnRngVf/mGvXwQn+VcEYysIXCrr+S3os2DWOBvsysGe7C4HSIu4Vd1tnWGHXGjrf7+1KG4CwXk+
3Qnc5GMwU7Ue+98wxZMlD1WO/2fLkMtg2Fb75qkVKuvqXW9fXVcTLpXWgo3JIFXfy12WHrwKBHFU
Dg55CqD+GU3OxZKgUYwt5CS26HXXDGzMi2xCp5bwIi8bkDm9P23pYJ4JIDSu3xvYcgAoUE4HIJGy
eBEp/LLdkoD6xyi8o5G7L577aPx9Ashk/Qpjvg7WgWN+ksWEZ8QD6thcQgBXzB/p6y34qDoeWGiE
FzFA0/vdBDuU9rGg2FCmesN8QdXqujg0si1doxfSB1zUskKuhACcEiXAUEDWBQ+ednqEqxUNwKwQ
dF2uuo0HY2eKC6hEE3Nq+Pzg+Gj2Q9TW4eF1eSsHG6UyEn4+hpZWMNjX7rQBkNZO8gL7bLDtwnUX
HUd4nLlxIgln2/RXaPSIETiZiPkUoCRVKY3r93ikeDKkyfgUGQ6YWI4I9gpXSeHYgCTsh7E2M6/o
l3IdHlW+lBWot9+8ysyBqpXGDKV3UtmXcg0ptq3iW5KHG7dN6q4xgUBswUyNbpszHu3X2EhsNkVY
/XcPsd+ysbI4A82oZG/A0MuCw7wnH15eVILVMjn0d5NwkkiQy5MSueH0f7I0kzOWtcRVMA5sRQ0r
eQtqZ9/93SqjbDrN6N6R3MVGLd989yVaKvcYPSI5yhIN0QiVzPI8VABiDQLpNWBEQYMJMNOnKf8l
WSOeRMGLWxua72YfIoKWojsX+cjH5j8a7o/AHtdj3k3Av2aNYdEBIqYnU8maiFOvMoXxPBELoTJ8
NguVuCTAxPCZn5IRgTKJPg3JspmZtsqSzbjm1iwgt1qFo1SyflQ7Wp0XD1oRbVIkTWT/j7Rj9BDc
c95D0tyN5RYewH6bhS8P3hBuXBMyv/24BubTa7e1nMvK5eqwLW7FIUXwL2vO2Vx5VDEuG09lVQqW
TlDC6yGw32DmsEsvgBlu//bb7DXtUH2dzdKFGl5kdlqsSyf5v9sAA9R5XZLIlTYimmhE56hg9jmp
Qy5dBSQqjJsgRH1LxCBKpET7NO6HloamkMgoMtMct+DzEhPb0cCCMMgl8z+Q53aGTqRJkkVhR+0l
99KkTpKZrMT+OqCVOpC1DoTpJVkKnpnffKfFCVZ135B/5Q05cKYGyGKF9/TCqV6RuutHCaJR9ZlF
OIjkbYO5AccOC3HiWa4o+z5CiLFDp2yIuNxgS9gnmmslUua7pf4ucPTLgb34fQbMoRT8whfAoOjl
W8wz1ADcFdfE82qY1g23R0Pu7XMGJEBuJoAs+Menxzfnfa7VH5+d6txE/Ck+QPTWqNs1Iu1ZM71o
87HHInRtXck89Xe/5kG+O1cd1joR9OBfrn98wbrlaqKf/c92mkBFjsmkuddfNsPB+nXNQ5McPkGK
hygtF5HH8QIso0NzXpFCWYq+tnpjAHFVD0S/ENq58F5LLN8Lr1FxA+UZ3xoGq6CXNIt+LTZ4SCF4
0gbfhgZZ47fstLoMfVgQi7SRbc3SHH+7FcauIbVIzTBT2hjNKts6mOJJdhK2FR30GVwbYuqIMoo8
vmonb2eTi6YNSTYe7/+dyA14r/okm+M0enkgSIb5bRysmDiGkn47Nz6bUauBBkl9gmQ3t57U3Icw
LZ66kBnvjZ1XhUpib19SNObjj6SRH4mGqWVmjUJbNQxR3+JAAl24mZbd75SwQx2JIpuIMBgL+h1M
rS2EnbVASrit0rubmFJhYV1zC/rjg224eNOYjEt4Emco7tdmu4pMy1vULv9kQza/v18hr8jDvEaA
0nUnF4lvb+IJt3jZWLMAXIcu5YWlGiyPbEbqYaOeNZIbjdp6pEq9J0u8H+Q8WXbI7Fe6S9xFEM/4
/Ab499l9t/8AjkV7LbS+IZN/Y4c9k4CJVaD6ZN0P+HIu7hig81o1ntoHK40rzo8oQ3HW5roYakcn
5dBkNBMoVvDbu7050RW/9W2fx+yg41pG/g5MVSVl9ANvR03RT/zcf0LScp6Gt050dtKu9jcVS6RQ
FdK9cHckRSKTP3eyuiVVuJ2bC7bmqUeOmo090AnNqtoN7HvbT/wfxzxUFFuFpSkaq11zeIGq9tBm
9bn+Mewkvv1HzC3qnU0xd2MtASHh0V1FJM0yh1fMK3dZHxXQzXA/pNcalcomDRA4rc9bMKohPiQ7
UEwc8ijGlq4gkwvsp19QLodEKviXgP5zsoEflAEb4Q1vt7+BT5tXa5M9Jr+ELeY4AZXgbIn7iZ+K
Sq8zjvZWTahUy4o4zw/mAxKLWtjXFqzfHIQMieK99uD4JAET7JrkNH0SEMibxqQP2WbbWf5Uhw8k
mM/ns2gpIa05jkO3MKGgwvC1pOzLr1mXOg+AKyWBBu79xV9NLpPFQ+M6eUIxmw5hOve9S+hgc5Gf
HOEcnBKdEB0ei37zQpAVQqFkUUmYS8vajJXfRm1KP2qKVBZ5w5Q4if2+FH0elLSF6SD9VgNKekRa
hJYCFrYA5tgffcenT4/58ZLfs5bbG2CQaXlxLZ0CwlmyVIuzZT79TRXWHOrug2t1L3adX63oNfCI
4/mu33qeb+JALXqCdY7WYRHUaY5ckfjAgfHTcR5Xx5T/RFuQDOHMCzKCJktg15s/gSN5+laXt42J
0qUhb2dezbxE/DeX131Q/mW2hKLMpj3tWSPkSmLrotWR1007PEgemJ10fyYsv71i7gXgEkxPAyHY
iTe1wtc4J1WDiqRlZE8xcyGvolQbuEAl+cL6jp8OSZHQSkTa07bgz6A9/PEQ6JsSmaZnaFslCy+Q
52felGCsZ119V41jfFwV+JbWfFo2HMQ35YT3maODY/ggQViCD55sPkJ+E36g3iimktOPEEW6qDBE
imKTBWV0s9t739sARBN1f9JKRDh0/fi02QJFg/t8ZdLSqyPtv0NOfyRjULdntivE9628mu8nRcv9
GAVOVBlyM3/AZojua8x8zmRoM+jDq7b1f+Bb0vGED4ZdKmo2OKaPUQmL5K9cY8ueiCX3PV24tCor
dfY/U/BG1ZZePoJEv3Yh320VXd2gs8NRCCbLLvQGvAIQ6sI1Uod3MqoNeiSaVaJz2qA8q4vVc2aZ
QvTeaj6ofmUVcwKcpy0ygh4o4ba+bEwQsOsmJA/pnIFRa5zFzX0FcwhdkO9peubuxSm4f/2gmhaz
wOGsqMNFiAhRTw7G5RVf9OWVQK5wPaPLSDphDRbfOAZITPdqtTZshzCsBlWRMcbB+g89JZWC4iBw
HVnN/yGNll1/wSbDwi+4aurHBFjgQYflYZiOzRzq7DPH9QAeXicsv1mvu5wkyelytYzgeN0f5WvU
fsVdj839zkUWHoTWOYaqHEjS10vt+4FCQrm/spsBqwPgXAl5flO2zjTW5RvfWJcl2VzBYGm7H1g/
oHZ7TXY0DBwuUlz1MDEVHutkSVZLlJcxx33sN1whQYPQw1lPX+97oGZa0vDpHy+uBImUf6185bUM
VCFDeXiy6gEF3wvq8hg7GJGFu9M7pDjaX+UzGiqEgsqWu1GvhEDX1TUrhRoVJ3IA/9AYiq6lQxAl
iTW7WhvAmwj569/Qt7qR6j3e2/Wy0hY6q2eMEh8LNx7LdIiFVAeQ8gm7hy5psW/PLY9hV3Qy8LAb
tmiZJ+Ak3uFvR4Z5YEM+XjBZCbhAg7vEOLtLCI20YtAeXA6AwT8WyeQ1rawUK53ZwJ/56W1jH8bh
w5QdZBHx9JX/xFMKNwX3YhshmgKtuGQFX4pDeH7lLuBknKXr0oVAqloXq0uwX4vvf1CsuvRG5oOi
8tOcvPUpamsAMccaY9mKVOiLUhG9H1keVUUf+2CoY/h9FVw7sqQpCpeiWvvm984mFxoUlcBDiOUL
VI2P+/4GjbwYXJ4uqWYMsf7Ndgi3nxUdy/4Fxs7GoAJ+sBzbM3ZCtU9yMLruGk63SSRtX3/A/02L
+ir1Wuln2shWs9Bztp2MRSJyLyOJOZd/2RuJ9VWwN4Uy3U/VydWeqpYQmf1dyExTJqoWn/wigZcj
7tASp3pzb4cKfEtVCSOby4ObHcAecwoTWbkO0jPou0+opG7t5yzlpooX7+q8ZynVF5HRgE1SWkIQ
I7Q7MwTcrKBPJCsP9ZhsnUbzEW412sH9rvB5XNmYXhUAeVqxbX3DqgjPit4XETSDkehQaycnYg4J
YduZeiuyzGUflJgOiVnQYUTXNl8xFZf3ips1GiveTKu8BMQLlCbH1cMt/6A0y1znyFFBXcP1RI8s
XH39dfZxc/xRQrfNiivaTvwDALis2bE5eELksDFZxyQpi7joPPcAz76xTE01pBvTCHzzM35oG/vV
Tp/vFFXBjufsYgGd3d1Z2AkozVUKoso7OUR4Ij1UxIkaq9oZP9sW13ijNcef8yVq0LPR6qD7cEvy
P0L1IM33IFcae+XTr4u+Tyh2MPYdT41dx/oKagmjClrC6Rnxu/qS3uFqI3SScBTsPMnbPGeSX7IV
cfrYEGS6fQvZ8sIaD0mTNce9HnTGYIwC9ZbuXa//OD6lAvnEtR/3bLLvFSvkQLODp1gLOxrpKf6F
4ACE1TVYg0FbpZTpMcmM5bkqslcOYzo6Ivm9QryGDP2TFfbaPSAAYglGjWempwqrA4Yif38VDugt
qFGt8vMSXj5TdWx+giDHj25Et6VZ9XTaxFEpS8tt+TAz7IxlyU5bcXIcuvw7rfwfVMrO0QrGS99R
p9o52u0wInO4eTZBVGeEgQCs0zoDgAL+Fbki2oMgbaME+2UDkUVaG1M9pGYuA9o9UfY/fDzwUOgB
1OG/HOmk9AU+ZUdV6ZwBXI8K8CeDVv7wSRWG57Ut/U9b/3RYYxVFF9WtZHRCHWyq3Nk6ySL+TzKQ
snjkerizY0nuTrN//rktzSwk8mKtHBu2yPAhrs822Xcnv1RzJJ46JKrvhVBEJTMuvvOMegFWCKGo
vY5wivT2P4OHLejMnEK/C8kMjJ/pxzSy6gBf/jFQ+5DXEEFwx88rR4r2FAXDCJK+15B0xKZEm9QU
OATqDRayf4lIlzagS95k5cJHQ23YYWSkF5IpA9QDtgTiXlLdQFz47UdtW1OqqwYRFooAoFndaZGg
koz9M3oBNH5XZo6Fb8MPFEtdtkHBXgxbkjM799sogHk15sJwRrUwxpMM1vx46wVyUjDFas/SuNgX
uwltaAQ9gOg5BUiTu65Lv4WnDKWvhXi+TgIk2a+3QuGI5JB5d/HS8b/xYjampvoKZFxZaLbHsPhe
I+Zr5JjPUBvUL9t0RdS6f/59X91mUH/XO4Wd/kA8KM3dw6k5uM+SCegOWDTl53QZ6V7olc6xoa1N
wRCrdjWloci4faqvi+qL4BCQBljLnzls6EbUmB1aBKpreBX+zTeg34svLD+kLSmwHpz9CfNc3iub
Pp18U0j/ZvRNHmLV1Xx4jfv/+VSZAeLJVHdbAj3O4w/fLdY/LERUEuwHpNA2UgzyhUhYu2vBPZtW
ZBeD8jRSsa/jwVd/Zm55uN9qtm0C+j2fhhJa+rqz6x3sNWUFeBCrZKkCEqVXTUzATixIGk/u1jcm
cYGCxBM6FFnmoXIX4Q6MBZzx/ICnNVRGM61wFqvWZW6wl6eSTyO5moMI26JTtKk8TExlE7Hx15GD
wNYLyi/lFokzkuQTnyfzICVOlxYi7l6sEVmfAS2+Dzv3IeEVPEskdKp3BQTeD4mxG4Rl5wJZm1ZJ
wO0vtF8Q9UbNBZuPOqlBvsGvgujZsqAkDpluc1FpiDqSE8SF4M30VIRTXQbG4ZmgUe/11SWrp5DN
Ve1mpEP+7dXJ4iQgvuXs7A6e0NEPu3ETjhvBxGlBjrndwtshE5WEE8BXcnggh8eW0i6leZ1gwmdl
58O09qlptxGttXt1r0MoTg3jddV0PGxNFbybJ3KRs/t+Wo7A//9Bv4VYSk/gakfrzwJ6a5yEv4Pr
S35vQplO/7jSNUVpLfuPm1TA2fLwRFug98YkE3diohJeCqEewhdMxde3DHlgbtca143xZGv/TEVN
kAGdK+SPcKfT7HvaIVds4IBD1WB2RpNrQzhpxpSX0rwTloHVotuZKoJW7Yb+H14IjNcBR16Ov90p
W9yyciAdWdGOTykFVCKKqFn2y3fQe0rhBzpyUMUabwPKfm2flH2zuwZ/2zP6Y3WW40Dq7iPcGrmM
3vfMu3UxkbDH2aGwTvu0l5hI5F9o3WaF885R2OSr/Y9EuoapdQQ6XreUZHvIUKBHOoVB8Pdrz5er
Q//j2oDL+BNjE0iAujbWcBANtX/xPhEgGIbNSmxNnnu/Kog5SX/jZ7CjCiojSNb8yvnUpoVy955C
4z2UnCyWC6Ma5xbm9PhKZkbqIPONaEaMBBDRIKBkAQJbrfy8oIKS0CX70FH5nZteg9LoSAUhilf4
XsrcgVNY5HZpO3RvPIXu/fTISDRh81AV2GP34Pd+kXrD8gcwWnCGt0NkiANY//JgrQxdMfPNWLpe
9jAVQU7mR/Mpp2UknliGn6r/DyL575Ey9XDhJB0eR9cZZxJX6IqlLc5X/mrSdcvXCsI3IGKdDF6J
y5P1CWwXRdnJKCVNZcdDSYyXhq2WU3eYONwP9MF/27HtP8vidkNc88MfwI+fZGhFSfgf86qevIOs
TfILo8Z0OVdJNTsuUhPJg5FngV4QGcrXrxzj7XybnvtgEHBYOPIyB8dCj2hjt08gsQddyRD1H1Qa
jg+qqmk5lFjw06EtqGJnStpRcC4+HUnv9vRi7Lulgjzbl8DSaVxOzG7rp2xsWBEpeqsQvNcSs/a1
o5p95EONrvCrPRUWTsDMimGaA+/YNJhA46JrGhwtIIycQ+IuZtu09Gt22hZTwDDQgIwb1xWwaTNr
vdwNekOl89tSTGWKj8+Xqw15hJdLv2u0doq6tMGKu6/HHRobHXRpNVHgGkXuvNgblraHW80TsKgL
RjActuUndWQV8aXC40LVM6CKMwaknXBmTqxd+vMzTAW0jT4sKHQUBQQfaHCEyNcWW7TsHxqbYG2U
j0GjwJbLZqV9Dk32ReFkxxl1GNLRZJ+1Ar3jTQ8pS0kniM0wdKjIrXTX1U5bzS3lCMmLryYFsnNb
hDpCuGYpyKjVtgLeTvuJ0cMLTVDkCOLncws28Tv7bJGVMl9z9IKtJGTM3yYOgCrhmqedb3bZ4JkI
fd1Ukiyb0PXgDQLkKP+c4h9Ih509TQBXHqpR5KcFO4Js7GzsjRQdFI5xbJyEVZLQna8qzN6+hZW0
sZMsOiJ/wn/WEmMoYgaXkX6d2pplVt6MIws29KQeioU3Rp7Bcjwb+1QN4PAjLxsJZUkZBDbnVuth
7Wh5AZxUolBDbtUE/P+IEZBIb3vyN4ctj390yAU3EAa9Z05i/sFnO9LNKJDHqJC9VQtf63uZA1Cq
9WNA4DeXDz7go4ya6EvlHkMBhoHVcXoa1JUPTqRthMOxA19vymgTkfvo9MppFzPJxum9eMDy2qDg
bmw/Qf+K7ai/vc/lzTsyVNhdpsDZOdPpqbAodEDYlV9NWHwMEk1alIy3AV2ACkh75nf2bLDr6am2
QfDOnOBv0DfXfqfbaXzZF9X7eB/EN9LSFXLXtoz7sFAmkihpAQQcFMo1NmxYvE1HLMmirQhpBPdU
/eh2d/IwFtXdgc+wA5gzd/v2dpBGEMFfRKJyQmbq4zetBewivN2YQ+eGMUUEsQcdORZj18r4HWc9
u1CcXSWGwfQSc7La05Gkr63S7JY4umS0E/E+eHB0nFy/wNa1q/6cWeaKnbG0waVyscLnErNdLETV
CvkCFoI4PoSRrosQhcU4cLhQWYuNL4C23TAzlhk9sInhNacmzZchg2sohAbT/Fx/PzSylvpmAADG
JpPiOrqsMnt9Ls1yCLc/Sf23qqdQkBzU3TDaczsPIEvSgz6dpSC8+wHyGHcJ7uVFRHLlJOzUHevR
MfGW9xQnXZ7Oyb0yZJgS+VMGlaiwOeqOAI2p6AW60SYauqlhHiB6CKoXwDxT+9ZWpP9AITewTEeJ
CRia3JOP1lNKk1LusEWSMyJR31IhjaLUzkpYHVhWcOYP7ukHso7GrZQPc+Q1VcCvAiG3I/C/DxJf
CJ5uPFxXnax+ssFzDlzm6VuaftK/fMnB/TAbwv7Fl4tx2350r2bxp93EoUAAH92OTmiDH4tcdoLA
/097jzbq+qNOSyeid0as+OdtLNRKscIV9+OqSsXNMH39ivQrXBPEKPgTDzqHxixTOV/88RPu0UgR
nzvlhKfFnx5BDcvsAKT3qyr0yloyKgXpl8Mum6Xw1fINHkoM0x5oDXwDBYokwcw8NS7cNBzw0WEp
23yrke35lSrN0DeDO8iEpj55mFOD7uYyL3CXkfWdIike5WL0xVM9J/HNUovVquV6mcvcPDgX/ipN
nMypOpCQRcQzDg/IaFB8PRf2tvMXmaEm945NNboShUdWtTI+ENA43hLxax3BYvAPTlfB/gFXdeYJ
goPEVyBzfWnkbDi62aL1avb1yxencX/DhWH6V6Cf3Jaa66SqJ0NK0zr3cUSLmHZ/V6EHoYceJaSI
E/epcdSaJRDMqomF1PyRy7eamFOnW1b3IoOkExnMTkXx1zWOCRInHO5GcnkTTyboYFgimrnB8AyW
eSaAJzWRZR9HzMKpP4g4qz2riZgnGZpdFxsK0iGHWwrlc6BZk3O1IjPFyhN2WhxtpCTE8jQiZfpr
aFwaNIej7UR4YSWcqUlIQ+2PYWQOS2EFVgkko79ejeHrkM39pd9uJdX5g8k8E1SPI3EvBcAIZpis
e1LOTHnomLXVADMwqeSWY8z13VuyNySn5HrHOlcK2M+Tih9SdN5+wHO/O8oD73M2Muat0ugz63t4
fLajuZWJEcgWm6D4ZRhQygZDxMbhiqlc/FFGQxhTZXoM0FBZGsrTUmZFNYbwBvu7r1Tkhe8/apfn
iGZgycetiSgPpDA9fvcSBJrCMQt29+bDE4WPOlmZE3vck3K519BtPOPEXTZ+3MiE1BVjFW6r6bxd
JEE37FCEw/toZOT0yz22p78snrym5WiKevBQRHDL1EbkkvOdXkqhAfkQuzgr40U/uCytPBlTFVVN
VTOCLqH4qDlHDSBBp3Sf2tSvVePahnNvlOyjWJSXn5MhJQEeC9vKu4VHk2tjCyVg5a79P+/hMjw6
lgELvoJFEOznBvv8GSqRti83wgzcxdr/+4WIb3Kq2AfdUpbVkRMVqnygxC1EVxOR4Xi+j9wBixx2
N483xIrVTIOZBfQZ+y7kf7kenTj4B0+EW0iMOiW3zHYvLsa51KSG7IDRGr4DcxX2AEXft1+gd8k1
qH4sd/VF1iEzGj6bVOM/K+PmcBOh4AFhZrhqgjHbEy0rYn0z38buOwkxGnC9dXe4YkOBM5TE28wP
SMe/ZJloJETYp5GEimQ+QjBW2OqtanAmA28WXtxKYgC2itCqTppTowFjm2fI253GYmJzGIziywSa
D3BJ0OX5gVijD/EJVC908jX5L1A6yB5Y2FD1ihwh/CvsPzslscky30fmo10pfgSjmOktlxfhbSSz
UJ6iAtYnLVDxG/vQOhmXdYvYMt/Oy+F8EIAouR9xsJoDeLxIcFgOkSFzTimojVTWUBxXX6O1bdBJ
hDKgYDC2ANYuUIZ0JCbZYPHwlIlsV0Yp6IEeEwiYl4wal5NZwdO9TsZTY1dAGMA6ByLtBIqMF5nA
+V+2lbFxdW5LcU+BOYrVJpZ69djhcf4xj2TmWHp6WL33WmJSQZVcPjkRumLdZQ83BYaXrloItMxa
q5lTsLaI1+fXW9Ybiy7wV2pOzW7bDJ/09OWEeeOQt8y4FjGjFYJd5uijffELYlSPN1PVVkLdvH5P
0RuZgRGhfE/3YZRnK1r6bOWKe1TAaqLInXMmgWzkFPVyHkVpKK86kY5ZZco2PTdkNA+Klo1Y80GE
4zAeE0iAtsyOE701p9o5OglDuTJlg1Jl9mLVvxtQsv8pcNQYJhu6frPf/f261Ohz68jLDPbalRPT
nZgcdPKx0q3sY1h4FCMjTSpomwX/3DuUeSptg3ECCG5XoVW0JDbfQIbczbjsiB5ehzFt5ZOn7Uf5
rA9hNb/XiVvajH2IjCRGHC/mdFyxtv8wl5GJ03p9W45vH2t/hBkxo8I3fMMn3Tfdt7zlatae8Xyd
zB0IQfP6lL9rOC+7/iY0vO6FuwOIDsYTrm2ZPGeOfHeHnxh+3MvndVbd+821nxz3RmR4arelpXcN
OQXSVLukgohxosHZGZWmU9RQrYvYW+Y6XWIBUVlgIOr8xDvII51AnG8xBkxcbG2v4Fu4rzk7Cqbp
1NQ0vVb+cwOXytdq57ttan0v3cL2hVA/OPeLV+oqY3PG0e26MeLTAJMAJqcsvGrB+PthTcTNL6Vn
oFsoGCSlg8QfYTfIxLMlO6M+1cUEYZZW6eauPMi1nZ6lV8gFOXZvMt0I2QL7+Q/fp3TTm/JVtlS8
70tK+ZlHhnNWJ8g9yFrvnomjOpnj+ICxf5UQCIewsr25BPHtQgRXAh4MRNANbY4+rIdK30GhNblw
d/e/l8/zeB2n2LAI1DvRM4OztMh8+hTjq9RweF6ayL3y4WMi89f8AnZU/YxLpUHUpur0JxWpwNWU
HHk+Or3RGxat+ROVcgAXjKGJQMnCNioTdHjnR/9Fn87D430i6z/nfARijnswNrvHrqArnL7k+ZaM
Zzv52V+VAz/4AE+7US8UWYTXkM0rDilMt62oy47hGGCw5tup0cIXjU7bbvGDGQHUB53sAi+d1LwZ
z7/07oEy6HiJUlowtpV/IzT0+9aTm2UeRcRNaQKp2UMB/dbf8ovTfsrsTC+pvyPY7R7vHECLKjfG
9jbDzWeUzJYS+wpERlLh+0mtJccwTq8T4n/gLmjL6hpZtPP5+B3PSv6mPsAeWLnzcCQOWuKPPoQX
c1uMyVMw7hay9OhzWZ19RWbVG9b8evVy1uzw0SNU413ULyBeEZs5Egbpt3tr4tHhCdmrvC0Hfp0E
WQkgOfF4A0IlhkuCylljAWGNsbO/0HKkY6cQWfwk/W6cKoKJ/fkl00ugTJBOOwdTgVMuIMW2C2BV
6x1vvr6TplDjeV62bKL365NTvUbmSxx7RUWx86LVA5K8oinwtIqmUmZ9kBxu8IhlU2Mb85g8c5XA
mEc4TJXz4gAW4+ptOw7sdydCNw133PVreQseoYqFIcXDn64hx1UAo4pBcQ5kXmSjT9veWUxIDIXi
eybAh4w0IkwYeRKYWTjVXpeLNhppbJXNDtgbeMzdOJ24zALhjLanvJtMqRNu0zu4AShqUVN/SQvZ
FX4EAdcS63GOBD8Fwgi/wicPoSDsYpe2qBliP1qn7AkEUAaCBrU6YSTHvzO/aMT2MO1hEM7H1IhQ
Ud9umWLITaEdtoRzIlpROoSOcZrpKFxcoLKBeAGF6TS4Tgm/9wtCymjLjPMMsFQVG7X+hqf98gx5
/nvIJW3+6LCNvJQ+Vd8X6lW4i8M3fSnv+iegh3Ztq7jMKWSBEKNWi/SFMJYHIPqw+mzY1QZSFPmD
oCXiQbktLfRuNdsB8ke/vz4jem+gdynpjmMB8jhyxoiXVaQt+EYw8Xmrr5bNoaRBeyhtG1wJ0xNR
zgLkbYE6GfI8EKOcczOvSzEqTMOxHm2bp3SjSJKIeBQoU07s7DvretUZMUsZDxINlSsgBYIsljts
BiUAbIX1HEuN2icQy5cHlF/BxK/HsbDpzmLf6TPqs1ZG5GBaRuiocS1gvwQxjnVgXQc/y8r/MISu
+VsTol0ewGJ93gxT946kMmtdR2eauGUp+EyHwfBAWnOVSHY83xiq5wcyO43NRX1EmTrp2hF2o//K
RAIn6FY9Nd/hH9WL9s/oiDsZcLx8smCCR90mcH8qbWnMX00hq/XLCIMPW31/QUMnS4akdOYSPAB1
qlXdgpKjgPb75H+k02Aex0oYGaDlHUXQujlV9IUdhSOC5uNFeKvRMm6zk6ZgS0QRATN0xmkYy+A4
Bf8SySxsOpWescOZyyaAJgwW8MSRxpBdJPnDoFh5t7+Q5BVlrvzeFo7EdKe8oMn3PYmo5MuMuwhb
fRYYR+fiDo06jeL3ZaFxOnLd84vue5dr1xP1N5lVAU82P9JK2ugThfzN7W2G44D4X08j5R8f7N7G
qROZZ0aRk2njqlEkVcG/CS/SZTPvCtMa1pNShS/h/u9p6C4wIL1iBoThTCY6DERNZ6AcCslyzU3M
bqjGxcZXNLYaaZtx8Qzx/drb0LM0Wu9dMz1m4lOvGLx/EfcEZ9nJ50Uyp0Lxq71y8B5mr9dCe3la
G4YUgRylNQl4VVASP1n3Vuo3AXZ9kvce2HfT6G9S3OdxXKBsB05ZGvDQHoj7d6uk5Y5QZ1R7zegC
9+Sd3OscqGoa+IO+/ctY3qK7AW60JoOvalLORDyy9jaOK+uVlvgeZi9YUFX5Cjrqpva00Pe4PxY7
aVWBY55OqbkqpKTi5hYC20UFuYfP2xUcldB197L771xNzTM9v+xmmxcP9R1nShracmoZnvVbnwC+
aoSwNXceTlmpl05kPyakn6h99JAUCgHUyGUZn4xmDwnxn4y4oOJl18w4eAeXSMKkJPwZsDlhw7xO
ksDeC8XiSsuDxOloN5muNwC03D3bi5a6lHq+6eE+bDdpliMPgzj8JMqJ6SZoCLBAXDFEVXy5Jo49
eO8yD7tu6L/qOBbU97nC+0xkjImPyxpOIB76+idHFvjnS4gZFKM9NXrCJf87c0f0uUvB62ZhbbQn
E0NSIcSWki5eBsKzl2acHVsPCORJFtI4MCKL8AT0KgClfSs0w61whM8BGoo2wvUHhoYJnHHHMBXc
lWHjXqFNuqcZYk9TwKfjU7ZlREye6zW380Cd8emVsbrjQ18kxqLUBYmw8+W4bGLFqrOLFOMfsPty
EPEpjT27Jz/ZudlFaUPkCHQqMV6K7mtOw/hm5BApOFh8AsTSMkuOSEksnsBGR/ZcwGIVz0wVPUe5
+yD9H7Ztkx5lx297OG1AU4Nekkz9U22hRv9t6UWvEeixPTXDt4QzaOB9g9UreSx5NslAAMA76ywV
VETB3H2ORspdvz/JvZcNRnOPe3E7d4iD7hBR7PF+7/ezuT507ajBPTBMTH/ekeOioURIb+cDuEH5
AzlN1rWFqam6EKNOZzCm4VP1QHyuIXpFOZbOTn8yCnaMib/YqAnQvjDNcx60z7ZCCAidDd256ekU
af5zo59gVgAwqqsZAM8lWLDjzb8/XntPRY+JOnwRjhsmjSlnHdlKhQJGlSScEEa/cB92lxKq3nDI
nNkC/Bflqy+kaC9sksFtMjg1detWec+EpkF3FGWA44rACDjuX3meAU/zql26of7/qi0ahfK1MQ9g
mKjRemntEw0nlGLlbhsAQYbumaSCwILqrONoS+yzPSip5YERBNUw/ZvWwWdxEaLVDHPFer3Ao89n
TWL4JxtEf8zoWQHbws6ampqLnOFhuIyVFJfPWIBBI5NLviF7UamCKkwfwmplvzSnFN7IE4SBbuAK
o1CEf2iYd8Mx1zeUu+/pjU0OW+8O+Pdub6brpEJVqPUpiidUjpGen+uQdcK1HpEyKyGTl0fCWn+n
SZoVDM1wcNEFAuT94Z9DbCHQL05p769mHNTPFf8iLEY1R2FexFg+NdxXLgy3JdGfdPpbzRZTGr6H
S98JWAHjd4+WXOdl+F3AiYeGdnhb8ovImTiiYZmy5bRUvg5CyyHAgnOkqFLZsPNU0Hivcbxk3h6Q
00vDBSvKStsHhJxd1zNgNKxHIeMocCalUQVhX+OKemeDXigQGDnwnNXjYTaTsw8cYZrEvx7JC2Sw
dPxKKbqOEQpZVPaaSdp9/BeHfm5IdP+clp+FzlFwPYWsLK89npjmsvSAbyEcxjl3OIRFhjkKWf4U
++gdfKX7oiEpvSO4e0cq8rGHrVcpvReZOii8sJhQvmbuDKQaUW8L/L4eBM0XH/mnamDGZsvLGMOP
nqQ8dYdS67vocqHphLeo0dUYxeFjR8iRC79zkhSmqlljiem9kOfQZjkO5y6SbH+9klNGM4ztxAG5
cxa06nQOkle07M9JamUtIfQ5CLYbzOq/qQxzq7Xx7UXgiud7S18xFXw7UgmSHf6u5F7MTPFWnqWi
ol/kSM9isTtqiQyklKHFbVMTLS1jQrTfEskAYKYW0U7Zq8AnAKc4Cuzx9qElD4EBed2GWj7Ia43V
p/TPUvOe1Xd/vcB5wQZmO7OdjPsmn5M9dxp2+/bYm/Va4EiTfIX/AYzUVylLKDCjOcLYhrkNDttb
vRXWjc7fx0oQP0cg2Wlptdk7yHp3tetc3OwSBa4BqveCBv52G9RXBHC15DPKrqjIcVWAS1mWFL0I
/3QrvLJJCBXkRe6dPqgaqmU9vIsRHEhzfkqGkyHrbV8F/XUvutOSnZWl5LyrUJBB+dZNgK+FXo4q
M1zBgm6RvHX2mLcuYE7FZ9726EOK4OQ5hRa4lGKxB6YM7oDFZcbp66UwHd3lFJwbZgUAgfhSl7gv
oX5C3cF9dJCWKcULNeF0o2zfiShFqS9VKgltGET5L+2icTlGVxuM0ap9MLO/gobx06Ib+uwQDT7w
2dZI/lK7TI03FUYKvdTBsVvYTmAAGPoYdbZYfiIOkOgD2fZKa3mzjiy1n/2chyK0cPpgfBGJAoxP
BDH37qdftY3xBUNBkTwuQcK+dmbfk7kncb0RKyP4RMSk/0NhwJ8qN9hbRE9/M8Wpxnu4NuG9T6Gf
GBxQLOabYS28PxB5sQP1QPpJUfN2TiDuwr8QYwXccTc6nA+wra3H0GjES2awcyVfSh2du8h03pyh
Ab59v9+7ilB0BkOCx+OwzYwMMNUArTO9anRi2xE/6sAbet8vEczvMYMY0WHsy2drPkaWNuOQmpFA
2jCOxbV6Fytwg+WhRyiIKtERMIgEomOnIaq6mqlUWkruaYU8RFclCpXiPTbLeJ0xFju5LF2PxUeQ
45EOzTXRiayU5Uwjp6BCfMS5kezCyKV76lXHaxZt/8msQb84+WKqcsiulT/oML+Wia0DZaeBLY5J
eAhixuFSmnOvzaHQQEfWpJlSKcYODmUXGAv54/WRsYEZ2VWCM2eBWggW/BQ52nV/2oc6kaL9NhDn
H5lTFx2e5aWSykFwdjtqxO/CwFb0BRXXp35mfZ6w5Nz0UnWtWDCxhSsOx2NBe6MAaN7SY9Q9PKDL
+v3LJAyrFMEmmswJJZWaxgrIfL4qhG6R9U+LvuUlwj/+g8MgZKGuDbG8MI5zmkDGxaHxzTwDoI/V
VrC9T3FyAiXgNXtndYyIW4xenwGGMtug5eojeTo7Z6QxPa1N5fGxTyo+BBxZa3qI1XUt9GQM2ZR9
CnnfnCqt5d4BhLtZyuLW5DHGh5CutQJvo6D7H6TiBEtqhEepLLXyBL6M1CDnT4fcd3uNxjXyUqZc
YKRgNJ0mJ7EI/p16YcjVKsQc+X4/2T943bgj1zKF8K/lukRphPbVQYZRNVrdsm/2LAYipy7fpbq6
1xUISrjcQbUvc2EO3gn85jeu6tvEuDIscrnykj6ugySUbRmQQLWPorTrthuMO+4DfsjsCK0n3UDk
OehGjKMHHZf+7tTPitREHty30N357375+BR8YYMN7sES6aGXGcASwbSUHtUg5FvmEu4dLfsCS4wc
qao2fR02VwQvevixRySQRbELxXIi4Va1GvAcPESOwgLlgaT7UvDG7fj6co7sGktJ1EjHaWFbjWcB
o/sUEQII+1HGmNKl0xBVnL4mo00eDkHoBM9hctGK4V308ZG5G3U2Q6c9ixMi/ov2uHZ13QaUhyjs
Nyq9vc4un/IXB6hioYWg4b0X4lNGzYSf7N4snlFOcAyj6NWmrJJRH1zYc2AB3nbglM9uJiCOv0Ep
g6FfKdWjsdGDy4XU7G8+ZnAGP0lQMuIor8l+0SN5DC+2iGbYb10Wz1ETjrsvhnCNsDFVp/5aJ2TZ
zPYoWdOuzov0vcnyZ44AeecmTbkt/wb2O4ZRwPXzLO0SegP8T9m0NnwVVBef3aU8RjSICQOHqcta
5vJ8V2P9o+sLnGQvu64VqxlCUaRZunCGYJFEu7YuXEq2N6be0zwHwhMS0gSvoI7seRGWeUr/seYI
/Yw+U4sOl4Oz/dj2/cncsSD5P4gt2q4HLrVtIdlYWB7xzuilZad4hp0vUyXIGk0m4PhI8aIHlPHN
EQkprp+CC0ZI5uZK7GTTEUlqnYkazZ/OYeqYIwLYVXxRS9+N+Ndcdifx87OO4mz3WNNwXPm6+wR6
mR4C56s5qEdOoMTeCepaiMQSVN7TZKJJf0Nur3XjPvde0MdhHlTUTkQk3hma7U8W257bOo0ni9Z+
rTNQju+HOuIKuBBGbHyB6XIxSp6efxHqmAx3/Httl4G6npvDs29qdmkzYOWgBYCP3mSdWyJpMpcc
jAgrHGkCdOMgHFWAxEr4VoRXjL+o7OLTQmK8AAc0uqcoL8iuGBmOhBGjGj52LWh8UWAGrEyncQBL
ZlG6kmzoEwmJObeEyO768fwwG/E752tXkRb0fvqO579gTveNRBBdVX/6WxQJb9BctiFYqyn1FVTk
TAvOY181jSC8NG8RXntw5nlwO2RMZAfPD49rrGW20o/7UueIyECwVWMqmWQtnNHpCmIIXuK1eOEf
XWXyz+5IyYffro3nhPbPrqBG1lsBd4PLZJ5NyUdXoZvZ7cEWs5O9IODIZXbvCAzRc2xdIf3w+web
1ZSJmREKlT+upBbyfEaCBghYlVFm+6WPzMDRxhkLziXH4zFq+UnXLiMHimjJIElvrVX6xYRqnxmM
qpUzAZ+TpSNnMwHl/BKx47ItG9fDeUm+ios5vPt7bA8iRePa1cAkFh/4Utp6B9dQG0qnXgY7/UFf
3utfllG8uk2P420k+TAy+jX34RoaIaHLPPU01kSpSiG1gt3UOsLoO9nmqxB49SFoLwdc+3DH3vS4
oL3iLd1KPJ2eT/FQJRM7WWqC3G4CYhv+swViF4pHtyYT9S3Rov3L/QoyDXnFc9eRxXcGKIUSWTTm
j+WfA/PuDdn5Njw76g0nbtTgMZXkNb52iTAP5fsKfl+KmCqeVCUbvnDamcY+kP+qjbxIInHYp+VI
vpqTgnulGDoFQLC5vBdraqJrT1y6h0kxEKEc/MzmI5fWSieJ/7Ugr5njDa79/y4hhHXHU/aWdsFk
bblFBufuRQ5u14pUm6Tafdvve9gfdFZKBRQumPwMB0UZCN8OfQsVA9xrd+U0NX3ZEj1q61KuKaxE
mEzgnrMMnA4bsYUTZI6349AA/6gNnYfdlIgqtDBATJi4CWpTEARMy/qSOqJN4vvMjh+9PZ6FU3oc
fGXkXPLvtuiAolTt4zOXhUC4sXGZMW9XvLuvNZwZn2hkj7WIFvcv8PF/9L4ZEPmo9Y8pu4FvDHXi
aECUo9jG3Vca2Zq+lJ+v3JK1l4nP0aryhy033xGj0TGJT3ZxOAyvlHbGFZH5viCDQsNNBXVoda3o
ZXEWLTiDU2c3o6FOmnm9sU2F9sYrMUOCp5CPUvbZlUM1UYvHgL69WqAAwqLDIVw/KzioAFSZSwsB
ekB08Nf20I6nUwtVvU1DAOc22/zgD14J09C21eeBzEfDdci5/Mb2Yabh3yGiSI90fhkdA9th+O6t
koq0mt+u4YVyZ5citPBGaL5ug/+Es9GcfW4d2vqcKixuCoYyaEnyw+XDDuD+Rrwt2z9T3/g9MKcH
gBuhwrPW1+96ZXp1aFVjhUuPrysT9jz/Nzi/fXlsumx/IUl+QuIx01NQPBNVwduKpbD09NKSDvRH
ACk/KxPbvtv+eOvsnxb2HzMIPA78Pex8rOnZBRZLuTN2XJ5WCC1GPYnGkz+zN51sesVB6uoWpTtq
0YIuPsFrteLXzMDFeTSPbnFf21eyqpnz8659/jTQ1TFluXr9Rb95hyE2IfZSCktthMOkPAU+vmLv
0oC0NwSqZK/vtYPtVkzcbWQJlgDRWxP6UC5sKJAGrpeEcgYUO1Ei3pcI6tFivgVW/Rx7EuV95I4z
+V9RQQDiQ6ejGZaNvrYyJkbR0KmwtPPuBuLSW/n0Jm8F9f4sxyKocPB66r9lTBqkcTJ41u3bxsdB
uBFnTF0QMb3sOMwMBjGc11crYzcUIgQosxTHHALn4xYWjR2SaBUyKCLoOmA3r9sXd+JHJhf21nCa
12MEjlze+2UGudILs3y191PKww3+dRzx/0nB3MQ0GT3sHoGZzGabRUk+4UEFQCIdF0hA+wcwQ3Fw
RLQwssbGfic0E4HmjbrWS5WLcteWV0F90PZO9+LAZOkP7V2tIDMiLLSoJN/8rjHfIRROgYnQ4y2f
b/mZicN34ajr1oZVAWpBQOKbrLVZL1denbKcE8wddn4uFByqKyusymrlqzr75U0zJJyqRvZzKiJV
hueuAQYPD1MCXta4nOFYB2U3fhsBOFRgJmjvuk7jhw/chU6BwMJegTAmYTOv6GIymGBa8xIrVfPi
E/hExqsgOZSxl3SAAVhb/gvXmux7SSGyffwkRQVUayxj3hDLv/KNy55bLWpbnNAY0QIGv0whbQTd
lQxVtTQm2yF0CfyYiMXTacIKef/Gqk5eLK3x9CzIpk4k+8VzldGhmI0A+Tb8Ew6xeOYcmdYXcdqY
kOtJi7AMUi9pnA6Sli9yl7wf8kEYBMLdNzxwzCiRTXwEZ4H7q0MhpF0GMBgM0dMJjjlI5cBrnkLJ
ZCZIVDfAjX8FUAX6dRejlJqIpk6OMZdmok4XqjJANGHq8hO38X6wXiz7O+y/I3+sVGXSSIafy3cj
/aAm28mnKAlxdSwz2nsrh8wxXt6X49R7+v9A66PthpJFy7qEWBM7Y2vFg2NmNHdlgzMaA4AgywyC
8Vq23ce9yXYyUFaVHZtj7QT9Slvc3riPgTrgDPEnfHyLDLq7fSEK2oBHBCuk9Z1Lb+1Odoh/9GWD
lwaxTFpVE2EfGyB9LijxPs1TgDkiOK3owRP6f20MLkDrUAvWjMs5ib6bmCkKvQSWDQ5R2g4ZKy0e
TpF9X+ejghCFM2rbkUrCBNBU8cm+1jrMqPBXNfjNG81rHRU7V8E/u+BFM/6kFq8YBrEFub4RZ8iK
0QJO9oEnJ28KoBGEXegq/pj63xxsENrpjmjpkZq3c4VQgG7/M00aeQVf27SDi9mIvgfPErRVp9ES
nQ6OEF3uue6f6nJT4zrCPlVFoZm3J5B12mnkgykUZNmMj93O4iBb7PsDWwTxyie/XrvuNdGnCMMv
q9aSaxWcz2CzPmvg+J9e6qEAUw/toOCScFby7MXFTMEkm0qH6/Y9byYOzx5Z6PBj8go9XopJJLer
aCo1j2PEf048xhPX2kPmfCND3MjimvKtM97ArQfaD1rJlA95bzc+YJ8miV0oSrF0G5OVosYaKRIl
pRg4HOlivwSQAEudd71nZiEpHuDE5HJ9dFz5nODeopxldLTIpujDZVoczRKg9MXpu5dZ/GFSd6oq
zzEs7ZWPS4nnRdlWN3BpveTqmAmrOfUi6xAoHbIYeVESl8YsTPkUpRcdqXK4duAsqKrv9+Mb7SSR
qVEiQ/o3v62jAD4NgoTlVEmHBS79XXUiC939Duj4Z0wBXxuDI2ZMXCleGn5gnXKLpPqpgRgCsobc
LFgccoNtJ9sZD/vGqPtrnNDwn/j2impg2uO9NAWdmtL4+n+sy8JxltsAXpbVCWCyWBIeHkQ9Do8C
ct+eytg+VPxauN6taOTVUk00qX+sD84H21XWccLuwBroHWUj3fTlSao7zh91CpyvwOshTvbmMb3N
wlZ6300W8/mRS0SBubaK37TO5mqnUf0LPtqV1iD7ZNNU1t9MXpAspKJhnsPg1vaDrDrH0zD/7L3m
6R2/BEcC3kQcwVtxfO26rlvFly8ZBFPvugRWMBif19NBMXJ92Rq5gizvPfJSwQBsZ12SzpAUFLyt
8mo/5/Kxz2zI+SjhciNQ/q/nwFJzU773zLu61XtkQHsnRRAyGyTgA3Yy8guRgOlvuM/nqi0H8sk2
z2+mhxXe0plKMYJ6Nluwa3aFlsjc33T8eTQ/VGsQ38YhhORx+i8uayniVx2ar8WgI6mTcXTIsPFJ
pPmVdIcM+y78QONAHOhkwU5qRQxn0en2zUcvi6U1/69+AmsHzg7mv4dOQsrlcuc24gVlSKTquGzM
OAUyCYDF5gk8KXFRSmaSAbXXuiq8Um3bwtBYOdnuvN738pijjHfiNJcAL5AWmhT3AI/ebbQ7eAyt
QwNP75FvCix0P2bIBPIzaddJuRG7UWbW+46hHJKhb4IbOpatgss67c0/6dmY1fiUVNwfRrMJD2dO
NDFJkPHLcGEHgczQ+p8hOj+X6LFSdwJMvuTGE1Dx/S0AwITJWo/WL4XYcV7KGTOVOab3iNFBbgjc
1JY1FtfxyqIVU4uXLcMa2m64vi71Hq/g1Gd6Ps61TsnhgNMHm6NQ2Z8oFSGvcVuzl1DotieWATaC
vQxcCnl1SlpHjta3gVAwHmAP9F2VPOhEWMvFwrThJkDK/zpF9dGhtLgdmW4tUCbOJJi+5NdADmtb
iIq0XwCEbovRZ0Ic0g/7udxmOb7BnI+l7omegicOU7QLCMVKrfZIt9a4XdCcmGiLXBkuqphJHfOZ
BQeA+h+iok8BuAktYqfTbZeMVKzH6iTUDVaYSUVOQF3AccjvXkqen890Cny5AxseyXYZL2yoI7HW
DWBoj36rb6db/H95q5U9z+AXhwJW8I6WQM/U7sLoIufiCycz9/XavpoqEI6Nj9Di+vjXsKMSi2/e
aIG/G1NynDd2/lExeJ89h5fgnn3V0cXLZpqFM+IK2BPv0BdrZX4SYaqdeDiiKctfjIW6Rn5xp3cq
LtBhwZPDG+iT/eTz8rtKqpIUq4syzHh4Hy2OwkmbmdQrTJ/mZjRy1Stk25arudM10eD2qanhDRNX
PuAXBkDh4FoCulWJPeGrj17/ECPFO5kjc9HeS+8YtlxCakAtjCyHebPrLg/LAU8tLkjPXHzES2j9
TFb4ZIVDu5j8ATWs/j6eIiPpglFomBgsreDcD0hh4QlSnNeilSlip95hc43J2rxZUHw0T1JR4l0+
TjvrKuJX2D7HZhNrQ8Fxev7H5M/jg6x3+RL35WIDylGw3atck+PRHeDqegzRfm5l0S7JWGS3e2MT
X9c32lCO32Edmt9lDYDFtr2ciYEfzSytUN2iC/k/tMEhEQfscRJIQYpyTkn1fQwmIBRBpzG99znE
WVEun/335r2mQd/KwrjCIPbfajlx3YyWUVRvfZRrEcP5e0tZy38BYZnoWINfVGGCJxAk3gYyKWrH
hmFM000Wf3MF8n/3FUvYwMHVvwqECWAKtLd4QHjgUJ7C8xTtOdoS43E+Kp204qk3i6tVimgmoW51
4h2Yqw5vBKcZXEzRbHkANemTccVOIT/aDLhk2qTA5BP4tlfR8laQYZU5rdAgT4F3iW5p6kNYbmHb
Dv9GW//CXWZ6oOv/pfRDs7VcH221hFNp5ofrKzIIdfCjkY8jN1wfonuu8w3NkmscRcSey4GUJ9Yx
Ai5elVbzN38tFT9qtxu81wX9MMew2yJIJh24gUqhjjL3qn/jQV3xRVPA00n0AdxOi8FB+Zf4toHD
5p8MuFEuwi/rNkSd0juh5dP1UbbogftSdTpMUQdMwGi1/i9HvAcbA2TMjQDdhpgw2ZlvHEdGug44
OiKGyUQRCTxZvb1n11RHn1nanKtRfJWWYb1kLyRjdLcEk9oqmN6WcisrP1LE/BeeNVfSWRkulUzT
ErlCZZhOUqEeoAQw7lm0edSNQ8DyNhcRFkF+KffvarX1LIUTcyFDXa03Nqza/ZEcb3SqNoMlKV9C
cwznJ6O6DcnjPqLl0+EzhJhhS9eGmfwUERKWiILIbUIMlSEMekyMQF1w4YvvCfdvmVMSD8xYmVjA
gagGKPK0p/06do3vyxV0X6Pus5dbIi0horl9azJ5Kl6V2VnmB3GKNNWdZtHNnrdBtCjlU+ICE2aq
Ou8oTsL/UdByVwmhvYETAaqO91Wur8paQcpLKfrXfdjuqXAA/Jt/9GIa5i7BKEpbk1vbxTOugL/v
LISHutCSXaDH+G5JIzP5NqXPK/+VXvoKZDzZZ7flMeB8RrS+JSDMdrdgiZSuQvSgq+5nrUzrDcbz
l3YVDdmJy6VHj8TecceeV/c2p1aGW/H553rMx2L+wRs8/KdW3S0tKiwlj2XfeZw8T356yIm/0Atd
NQiuBvrOjmsDuPYjxPi98pACGnDWzUeDQoKhTMAIGZEiy4o8nxNlX/VKBpXnAkPNW7PfRWsOE88I
65LZqwnFX5UXCehHMLWM8pmH0so65y6SCVu2y+twtzOSVQP9e4A1RXukD409qI3SO2GDNu+Fs0lA
Lv2NJw3/ni/0XqKKi6r6Stqiv9ZBmHFqyfsslYOPboOmWIC5k2OsRvYNIrCAQ4sBlYppW1EGpD1W
nrdX3PJ+m6U7ByFHaLEpZ0wp376gUDlOnYUh+E71qyEG68GjEv0mHzrQSv0vccCkyV6u27pnayDQ
7NDDqo8aERj7+x4ohDq2IN4FsAMWXgSCUp/+p662909phfjPM7JrHAa2aiWeBhr/wAOSJWZNX+6/
pZ0mIuIWc8QPXWsHWcU8aNfoBUSDXYBp8My0PyYgRUBYnYvwJG53xU4OmlYD6hlg9Oo82MItJUwD
vo2hPE2h9jGaukNA8GTecvUSy6jEp537s7zVyyPOpsjN2s2XqEtwzCyF5BO4jifsUUQI/3sPC+su
5Q6ubzQKb/zkoKrXR3kmI4EJ0LN1sXY42aliXST/vpTZYOH5vlv5OofXccc2FMBpo7TwtKNX/dJI
7R5osyBt4sGIIFHoxMbCHAG35I3N4I5NM5zYaHHkbvam9OltbMyVQuOD0CBFkBnFudA2miuUEaDF
hIn3cJyjyvGSg1ER6efIU5OpIEsQ5eMnqum9MYWV3vicXp02P99Zqjo2wwNYV48PAnuCGip+fxRd
BBE/pJMr1dVBGqURMEOGZu//sMuG4ZOkBoQkl2Ar1KtNXBorzRBKc9HqAlw4uBbX8t7ck4WUKWtu
cxB7QRySGOB+w+/qu18eUXvarKA1Nss3W5JTVdwgG36uuhN9o2VTbNu6P432S/l3tR/529Fk5f5U
3NMK/h14so7LTeAPa1kNO3TvmBWTVlc4qSJSMvFgBhwGZCOiEDZ0Yz8oChNs4fHU9/of6o0E4DFJ
i1WDT9JobxRP3vc31Y+Djmpi7Fbqi/5Ef2RmH6NBNCvJ2dqGiLzuiOAFoywhauN6OGdndDmzoDPM
bcMy4WOwatpxUJl6aAEFZW1hkDemsmgeQ34UVhnMWhfwCa2wjB79WVrIer/SEtE1chxnWsXt+Mtv
gqYuDjVKIbY2pXZr4ftfy3oFwCi5wRYy8149oy894sEhoANqCQFgX+T86rdhpZj06AsyNoG+ahto
FfJXWVNRP1s3IshSwEjtq8Vy7vHEnA0ZUm9nsv1wE2bc3D1w5MNl8XxIjbF9sa6HoLPlVQj3K5Nh
ABHGcWegwJXGgrFqZ43AePsfQhmt5WCrnSduglKLrgbv6d6kcvC1TP97Y7tOSfHO1ooBLowS8K3T
m4spwJQj8q+LQp3TBpnnbJrZMpsr4jTcMFf5RbxE8npFK63jwS1xKwoHmhU3BiniLN0Xx4XVmL49
7YVuCgu8RN81oUF2qr8FXEjwWNgHffCq+Tgj++aALj2rOLtT/YzawCkJmFKyK6iGloWRkeXBI8uC
hKMuNrj7mNP4u7mpd+VeWy6fcnkUakaoe5W2/bJHiPyTSHLyYA0G4ocLp1EZ2yJvzxRUbLznhC95
WrnFmy/W21mRTmbHeBFRgE/E7MZbBRZJ+OXwrYHfWWEQP/nKqljt/8oxXkmLLq1RxbDaFME+RZBM
oNvjAQyauQHQfAUSLS7cNiNY0W1/M1XEknpZP9/qeNW1mGWvHGxDoKPDm8KoFRkymewkBgqjrRDF
4Vvdv6RqlW7Td4rYCwo9CrtD66lgbrUBThNd2XxbbiYiuc9zoevWHKZHhwysNNPE4gvEqmm5bRXx
wlwoyaSsinfl/ydtJOicH2n+fDfe8kPFWGQeea/Do6obqaDNE5LPUDG/HmjxTmk97q9T6B+5vsSl
OgN+5OjD/NZIPq79t+IYK32QHb+ZDlMOuzPFWrYvIN2D+trkozN9Ect8iX1Tz1sT1YRNz56OG6h3
7oSnAujlVM08QwVmSS5NE238cjTZvdCrUO2OfyJvN+Hjz2yz7YwsPewyHs0gXvXOtSyikGILH9G3
WCCEAEjCuAUh0xCka1SqYyvXoGYDMSG/APThrnJFrXcIakC261fHzXc0ZClSWuAmebPtFT9oLEmj
6M0rdwRSuDonPm7evN9rMlAsTuXzw1X9omBuIY7HC4z4C7peGZJt7mol/uNIo3oEfOV2kdBGvWdh
FcFdXj01OxSpiOjIgwE2ljA6cSuN4ThKKU7wquFtf2jkLxLknJZEGFkeGlGI6A79l1cH6nz32M6Q
hV5STYsUhesBGOzAtf65Y3r3Xp8UaGiEafK5D3bq3N52QBIlFwu3iet7nXUVnCLGYaDAYMCh7oOW
IIUWHJSNYb1FFM9J9chTNDv6smyVJp9Z9RXr0DILGZlQbGy4OCVJNn7zOG07ZQ3fhgu+Da72Q2jx
XCsk+tqzwn7gqsINOFQTswqQWUCV9rgtO0mmP54jXy9PJ2TvH0RpjI3t81FApSVH+jM0HaL0LIpX
9zmv9p8T5uVDxWvYZOE1tcX89iZ70evD2/BFaB9rlreIhUh7DfkzE1y8E6yHPxyLtXmxq2Evrqa9
wJg52hGnj9aNAJp/2M6oJH42LFb+wHgZ4uXOtQVYXEIhVeGlL4XfGWZqaXUZK3lQWl4ks9rh+sTZ
/DKOrY253lgyGo31RmUVK7TnvRLUytmcZKfk1xxQl0D8UyfkR2/fRNU9BNv3/U9pESzaIPODc0J5
3uG6aTSJQItPErSybQTXCoAN7bvrNJpEuVO01l5r+4JT5AKOAIwlvnUO20ugMx7uxuimyYhYy28f
9QvaFD77Mu0l1ijiQ+Xwa77JctFvYAFJkuRS6zaTst34rSCbvwhpCUfsFhpXPVT7QRpRDL8uzL7P
C1B4L5hpHianlNBkO3DDAL5VIfZO+igHrOoPvuy7e4kMHrH10ijf2bQ29ZPJpbOYwTW+2uZhHJWY
ShP4HVDZ7HbMGjfI7n+mhLI/MXCx0TB7p0y6dWSXNRzgFuP4LcAs1RtbFS35Atl1AbAhETUemaAM
GiLKAKS3BYLLYsOjw6W5SxwSwNVBHPEkTeVGbT3c01lHu+aLafRS3xUZUX75PTD6No7wJSZiQ34O
XnQd/ZIauU3fmZBFoToIhl4r9jIFHCTwbNKmjQVHir2UDqRwKNw6KbMN+5wzo6QmySZrxLhsd4dv
SOE4LWe79c4TMV4sUv3NG/tOheSPq/KRHhqYnAQC2WyWvT1ROMS+VEvjL7JdqENPesc+CtEj4Ktw
CndM5OUjNrTbaj76n9hJK+e1/KJvi6t8dGoQS1yHfl3cRFN4zudJ7y15GV83O9PNby57X/5RKHDU
p81lDnBNj2EFskuZbRMOV2ymoObwUBEK7dzlMJCEi+jR4oe7LOXDBrgYONV562uwrxzDOjkVcYkt
RBVEf1tzLOdCMd40Z1pR3fnTm8v89Cn3pWRe5KY+GDaMAgg4zO3db3LBRQbceT46fYsCWj8FNTsw
tX7Knq/IGj6iIQJPoTfi1x6pMscCGsU8EHA9yzLVRljqASqS/qZoYE0y3UXuv2tZdVLrFlRHGkyE
XOq+7bHVHDBpYGHzU/Ody9bIRgHzspFeLcPNpjM9v7A5FXcFpkoZu3niAbyrNHjaxYYZKMj7xHXc
tYWPQHps+g8UsB3t50yP1QrvByztsW4sqFqXMnO3FPrDZIw8z0m9qwMcu+G0enjzZxz75RddgnBF
jqInFc03C3sEqUwdnmH1965NCqb+pdLcCbR131KBcqpHxGM39Oy3nZRz6deYJ3ijVCcmz9SIYtlQ
E/mT3gZYkLKf52er49sGAVIAuWE88P/WO7OCUK2hRm+dGXwGSs63NZ1ifnMaSiEdQFLqXvGY3wsL
Ey7QaLQ+34snlXCffCE9VQNsoEwJm1YokFi8aHROzPi5uOM6/xsE9VAf3pwJIoH17M7Nxz9Z61A3
LVapE1m3p+xHqkEKxyLfUymxg0ktrr5BXCShx+p4hydVyRg1OBpn+wfh1YzqeXL1oMtjP6fBiwBj
ZFBs9zeayvE6Uszil4chdRIsJxTXHtC3oAdAPPW9Fpw2aba0drkEswbXCVowCWLuK5ex7x6AtSxe
ygh9aS5A8AbovjwSib0+a7sdvxXOtR1LoSyjHHgs1aVPkdxSx5PfJXQqNjHNAme+d0ZhwdSI+VY2
12UsJVzvI5eklYx8OiTpqgOKRbpkq5Th+ljexNWRbrK/78pXMzYHZAvlpcOZ8ntUn85VCv6xhLsu
pgYRiFsF5FgfaPwImu9fMu94UvHxXMXxkDJeH1hGvmo1ozS34qveCqDvIg8EHD5C3VTH//7W+Ntd
6nOpxq3hq33p4QPYuLzZz1blOlY/T515lnXzQKJPdNDC+celkWLn7kHEq1tf2cIs3Q+PMVNg9a1V
JvUTcdZrjHp3n18r0Sxmmw8k4BMNVq8eKHlQdcmjaI6kTatAnIb0fGF6PNNt9DX2aQSXjRBTzCrB
AOUC3w6qwTRadNOTSq2L3BH/U2GyfgnL1ePbckp5HmMYcA6SnZcbH2Rq5QI7vqpyseWKxCZr+3vO
P39etVa+gw8kKHws9ZW2rmK7cDNf+WsojCyM8d/j3fpcc4vUXMGe8ofs1L7N2Y9pKZNdpR2LVT+6
qEkeilswjqTP8Wfci8BeJKr1j9HZNQm3/vHRXJxcl7NqKVhn8eOODGuGTxHYN/euxhl4lJXqx2JU
fmQ/4YzqJTnBf0twIcrxn+SBdsMFdB55G3MOUnHkkYBmOC/lPI+BPs0PxRo4gd86xLOmBHZ6AihV
0r74BYTPQk2RWxwdTwjtQwdBcIkYNs5bGyZpOp8lvDEAkGpP0Z+g8wFqTEVvKT8UMmA5JpI9RWFZ
UJ43vdT/5vsRlqeJcDnlfgxSq89A4wHddAv+E1s7BTwA/9DLPuyY0P3EiPYEirQqMf5hA29x68Me
+OLhiNJgXUku6jX3QDM1hkmqruHP7DjpwnAMtLmNcnnkVOeSh4Q0o87f6GQd6xDuBzkUtPxuVNOU
LMYuzXL2vzpS2yB5RiHYWmoBV7aAC/P/xnWtIesvh9XIWv2dCfVjM2QFVFx3DFpR/X3UvOBRb0+o
C6IRl+pF1Ch8amdtBP4OhZPrMJfQjGnBz2X+FfAUP5a5qhjQ4t6kMIMkvEqlHhRukGmBEW2h31EB
WLyUgyYGyxTm++nyAELvuhjSY/5W2NcKs8ocKgInYjg/1qfBGN1fbQtSQJfg3MIEhZPn/RDTi5m1
GMJVLlW8NAkv74bTP1Kt6o44Nsc49lc8kACQOfDbmveVKYBv89iwpAfeuRkgB42qTz3Bm/hl0zxR
NpfB2Pqf2IIRQdQqmmJeZS9693cc3jfhZy2ihMzV8z5crESQGmKUS0f0ZPIybXUoOHjc6YDKkJmn
G9UMJKEQEyWOk/lZQdtDi5daul5uRw71dH3DbRoid9JPhocqBg2lrmj86YxjWKmYlnqd4UI55t3T
ealccrioPgVATeR3duBFAoiE0MuZhcWuNbf3vAs34k/loz5+PBAMjm+mcGeD6HWP+QF0llDDzLlb
agEjHvKBOl5lWJLkLudJf6vG/QcDl54=
`pragma protect end_protected
